module tt_um_dlfloatmac (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire \MAC.a[0] ;
 wire \MAC.a[10] ;
 wire \MAC.a[11] ;
 wire \MAC.a[12] ;
 wire \MAC.a[13] ;
 wire \MAC.a[14] ;
 wire \MAC.a[15] ;
 wire \MAC.a[1] ;
 wire \MAC.a[2] ;
 wire \MAC.a[3] ;
 wire \MAC.a[4] ;
 wire \MAC.a[5] ;
 wire \MAC.a[6] ;
 wire \MAC.a[7] ;
 wire \MAC.a[8] ;
 wire \MAC.a[9] ;
 wire \MAC.add.a1[0] ;
 wire \MAC.add.a1[10] ;
 wire \MAC.add.a1[11] ;
 wire \MAC.add.a1[12] ;
 wire \MAC.add.a1[13] ;
 wire \MAC.add.a1[14] ;
 wire \MAC.add.a1[15] ;
 wire \MAC.add.a1[1] ;
 wire \MAC.add.a1[2] ;
 wire \MAC.add.a1[3] ;
 wire \MAC.add.a1[4] ;
 wire \MAC.add.a1[5] ;
 wire \MAC.add.a1[6] ;
 wire \MAC.add.a1[7] ;
 wire \MAC.add.a1[8] ;
 wire \MAC.add.a1[9] ;
 wire \MAC.add.b1[0] ;
 wire \MAC.add.b1[10] ;
 wire \MAC.add.b1[11] ;
 wire \MAC.add.b1[12] ;
 wire \MAC.add.b1[13] ;
 wire \MAC.add.b1[14] ;
 wire \MAC.add.b1[15] ;
 wire \MAC.add.b1[1] ;
 wire \MAC.add.b1[2] ;
 wire \MAC.add.b1[3] ;
 wire \MAC.add.b1[4] ;
 wire \MAC.add.b1[5] ;
 wire \MAC.add.b1[6] ;
 wire \MAC.add.b1[7] ;
 wire \MAC.add.b1[8] ;
 wire \MAC.add.b1[9] ;
 wire \MAC.add.c_add[0] ;
 wire \MAC.add.c_add[10] ;
 wire \MAC.add.c_add[11] ;
 wire \MAC.add.c_add[12] ;
 wire \MAC.add.c_add[13] ;
 wire \MAC.add.c_add[14] ;
 wire \MAC.add.c_add[15] ;
 wire \MAC.add.c_add[1] ;
 wire \MAC.add.c_add[2] ;
 wire \MAC.add.c_add[3] ;
 wire \MAC.add.c_add[4] ;
 wire \MAC.add.c_add[5] ;
 wire \MAC.add.c_add[6] ;
 wire \MAC.add.c_add[7] ;
 wire \MAC.add.c_add[8] ;
 wire \MAC.add.c_add[9] ;
 wire \MAC.b[0] ;
 wire \MAC.b[10] ;
 wire \MAC.b[11] ;
 wire \MAC.b[12] ;
 wire \MAC.b[13] ;
 wire \MAC.b[14] ;
 wire \MAC.b[15] ;
 wire \MAC.b[1] ;
 wire \MAC.b[2] ;
 wire \MAC.b[3] ;
 wire \MAC.b[4] ;
 wire \MAC.b[5] ;
 wire \MAC.b[6] ;
 wire \MAC.b[7] ;
 wire \MAC.b[8] ;
 wire \MAC.b[9] ;
 wire \MAC.mul.c_mul1[0] ;
 wire \MAC.mul.c_mul1[10] ;
 wire \MAC.mul.c_mul1[11] ;
 wire \MAC.mul.c_mul1[12] ;
 wire \MAC.mul.c_mul1[13] ;
 wire \MAC.mul.c_mul1[14] ;
 wire \MAC.mul.c_mul1[15] ;
 wire \MAC.mul.c_mul1[1] ;
 wire \MAC.mul.c_mul1[2] ;
 wire \MAC.mul.c_mul1[3] ;
 wire \MAC.mul.c_mul1[4] ;
 wire \MAC.mul.c_mul1[5] ;
 wire \MAC.mul.c_mul1[6] ;
 wire \MAC.mul.c_mul1[7] ;
 wire \MAC.mul.c_mul1[8] ;
 wire \MAC.mul.c_mul1[9] ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire \wrap.state[0] ;
 wire \wrap.temp_data[0] ;
 wire \wrap.temp_data[10] ;
 wire \wrap.temp_data[11] ;
 wire \wrap.temp_data[12] ;
 wire \wrap.temp_data[13] ;
 wire \wrap.temp_data[14] ;
 wire \wrap.temp_data[15] ;
 wire \wrap.temp_data[1] ;
 wire \wrap.temp_data[2] ;
 wire \wrap.temp_data[3] ;
 wire \wrap.temp_data[4] ;
 wire \wrap.temp_data[5] ;
 wire \wrap.temp_data[6] ;
 wire \wrap.temp_data[7] ;
 wire \wrap.temp_data[8] ;
 wire \wrap.temp_data[9] ;
 wire \wrap2.state[0] ;
 wire clknet_0_clk;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;

 sky130_fd_sc_hd__inv_2 _1078_ (.A(net121),
    .Y(_0001_));
 sky130_fd_sc_hd__inv_2 _1079_ (.A(net40),
    .Y(_0000_));
 sky130_fd_sc_hd__inv_2 _1080_ (.A(\MAC.add.a1[12] ),
    .Y(_0317_));
 sky130_fd_sc_hd__inv_2 _1081_ (.A(\MAC.add.b1[9] ),
    .Y(_0318_));
 sky130_fd_sc_hd__inv_2 _1082_ (.A(\MAC.add.b1[0] ),
    .Y(_0319_));
 sky130_fd_sc_hd__inv_2 _1083_ (.A(\MAC.add.a1[0] ),
    .Y(_0320_));
 sky130_fd_sc_hd__inv_2 _1084_ (.A(\MAC.add.b1[4] ),
    .Y(_0321_));
 sky130_fd_sc_hd__inv_2 _1085_ (.A(\MAC.add.b1[5] ),
    .Y(_0322_));
 sky130_fd_sc_hd__inv_2 _1086_ (.A(\MAC.add.a1[5] ),
    .Y(_0323_));
 sky130_fd_sc_hd__inv_2 _1087_ (.A(\MAC.add.b1[6] ),
    .Y(_0324_));
 sky130_fd_sc_hd__inv_2 _1088_ (.A(\MAC.add.a1[7] ),
    .Y(_0325_));
 sky130_fd_sc_hd__inv_2 _1089_ (.A(\MAC.add.b1[8] ),
    .Y(_0326_));
 sky130_fd_sc_hd__inv_2 _1090_ (.A(\MAC.add.a1[8] ),
    .Y(_0327_));
 sky130_fd_sc_hd__inv_2 _1091_ (.A(net43),
    .Y(_0328_));
 sky130_fd_sc_hd__inv_2 _1092_ (.A(net66),
    .Y(_0329_));
 sky130_fd_sc_hd__and2_1 _1093_ (.A(net112),
    .B(net40),
    .X(_0002_));
 sky130_fd_sc_hd__and2_1 _1094_ (.A(net40),
    .B(net105),
    .X(_0009_));
 sky130_fd_sc_hd__and2_1 _1095_ (.A(net40),
    .B(net119),
    .X(_0010_));
 sky130_fd_sc_hd__and2_1 _1096_ (.A(net40),
    .B(net118),
    .X(_0011_));
 sky130_fd_sc_hd__and2_1 _1097_ (.A(net39),
    .B(net117),
    .X(_0012_));
 sky130_fd_sc_hd__and2_1 _1098_ (.A(net39),
    .B(net116),
    .X(_0013_));
 sky130_fd_sc_hd__and2_1 _1099_ (.A(net39),
    .B(net106),
    .X(_0014_));
 sky130_fd_sc_hd__and2_1 _1100_ (.A(net39),
    .B(net113),
    .X(_0015_));
 sky130_fd_sc_hd__and2_1 _1101_ (.A(net39),
    .B(net108),
    .X(_0016_));
 sky130_fd_sc_hd__and2_1 _1102_ (.A(net38),
    .B(net111),
    .X(_0017_));
 sky130_fd_sc_hd__and2_1 _1103_ (.A(net38),
    .B(net107),
    .X(_0003_));
 sky130_fd_sc_hd__and2_1 _1104_ (.A(net38),
    .B(net110),
    .X(_0004_));
 sky130_fd_sc_hd__and2_1 _1105_ (.A(net37),
    .B(net109),
    .X(_0005_));
 sky130_fd_sc_hd__and2_1 _1106_ (.A(net37),
    .B(net114),
    .X(_0006_));
 sky130_fd_sc_hd__and2_1 _1107_ (.A(net37),
    .B(net115),
    .X(_0007_));
 sky130_fd_sc_hd__and2_1 _1108_ (.A(net37),
    .B(net120),
    .X(_0008_));
 sky130_fd_sc_hd__and2_1 _1109_ (.A(net40),
    .B(net2),
    .X(_0018_));
 sky130_fd_sc_hd__and2_1 _1110_ (.A(net39),
    .B(net3),
    .X(_0025_));
 sky130_fd_sc_hd__and2_1 _1111_ (.A(net40),
    .B(net4),
    .X(_0026_));
 sky130_fd_sc_hd__and2_1 _1112_ (.A(net40),
    .B(net5),
    .X(_0027_));
 sky130_fd_sc_hd__and2_1 _1113_ (.A(net39),
    .B(net6),
    .X(_0028_));
 sky130_fd_sc_hd__and2_1 _1114_ (.A(net39),
    .B(net7),
    .X(_0029_));
 sky130_fd_sc_hd__and2_1 _1115_ (.A(net39),
    .B(net8),
    .X(_0030_));
 sky130_fd_sc_hd__and2_1 _1116_ (.A(net39),
    .B(net9),
    .X(_0031_));
 sky130_fd_sc_hd__and2_1 _1117_ (.A(net38),
    .B(net10),
    .X(_0032_));
 sky130_fd_sc_hd__and2_1 _1118_ (.A(net38),
    .B(net11),
    .X(_0033_));
 sky130_fd_sc_hd__and2_1 _1119_ (.A(net37),
    .B(net12),
    .X(_0019_));
 sky130_fd_sc_hd__and2_1 _1120_ (.A(net37),
    .B(net13),
    .X(_0020_));
 sky130_fd_sc_hd__and2_1 _1121_ (.A(net37),
    .B(net14),
    .X(_0021_));
 sky130_fd_sc_hd__and2_1 _1122_ (.A(net37),
    .B(net15),
    .X(_0022_));
 sky130_fd_sc_hd__and2_1 _1123_ (.A(net37),
    .B(net16),
    .X(_0023_));
 sky130_fd_sc_hd__and2_1 _1124_ (.A(net37),
    .B(net17),
    .X(_0024_));
 sky130_fd_sc_hd__nand2_1 _1125_ (.A(\MAC.add.a1[15] ),
    .B(\MAC.add.b1[15] ),
    .Y(_0330_));
 sky130_fd_sc_hd__or2_1 _1126_ (.A(\MAC.add.a1[15] ),
    .B(\MAC.add.b1[15] ),
    .X(_0331_));
 sky130_fd_sc_hd__and2_1 _1127_ (.A(_0330_),
    .B(_0331_),
    .X(_0332_));
 sky130_fd_sc_hd__nand2b_1 _1128_ (.A_N(\MAC.add.a1[14] ),
    .B(\MAC.add.b1[14] ),
    .Y(_0333_));
 sky130_fd_sc_hd__and2b_1 _1129_ (.A_N(\MAC.add.b1[14] ),
    .B(\MAC.add.a1[14] ),
    .X(_0334_));
 sky130_fd_sc_hd__nand2b_1 _1130_ (.A_N(\MAC.add.b1[14] ),
    .B(\MAC.add.a1[14] ),
    .Y(_0335_));
 sky130_fd_sc_hd__and2b_1 _1131_ (.A_N(\MAC.add.b1[13] ),
    .B(\MAC.add.a1[13] ),
    .X(_0336_));
 sky130_fd_sc_hd__nand2b_2 _1132_ (.A_N(\MAC.add.a1[13] ),
    .B(\MAC.add.b1[13] ),
    .Y(_0337_));
 sky130_fd_sc_hd__nor2_1 _1133_ (.A(_0317_),
    .B(\MAC.add.b1[12] ),
    .Y(_0338_));
 sky130_fd_sc_hd__and2b_1 _1134_ (.A_N(\MAC.add.a1[11] ),
    .B(\MAC.add.b1[11] ),
    .X(_0339_));
 sky130_fd_sc_hd__nand2b_1 _1135_ (.A_N(\MAC.add.a1[10] ),
    .B(\MAC.add.b1[10] ),
    .Y(_0340_));
 sky130_fd_sc_hd__and2b_1 _1136_ (.A_N(\MAC.add.b1[10] ),
    .B(\MAC.add.a1[10] ),
    .X(_0341_));
 sky130_fd_sc_hd__and2b_1 _1137_ (.A_N(\MAC.add.b1[9] ),
    .B(\MAC.add.a1[9] ),
    .X(_0342_));
 sky130_fd_sc_hd__nand2b_1 _1138_ (.A_N(\MAC.add.b1[11] ),
    .B(\MAC.add.a1[11] ),
    .Y(_0343_));
 sky130_fd_sc_hd__xor2_2 _1139_ (.A(\MAC.add.a1[11] ),
    .B(\MAC.add.b1[11] ),
    .X(_0344_));
 sky130_fd_sc_hd__a311o_1 _1140_ (.A1(\MAC.add.a1[9] ),
    .A2(_0318_),
    .A3(_0340_),
    .B1(_0341_),
    .C1(_0344_),
    .X(_0345_));
 sky130_fd_sc_hd__nand2b_1 _1141_ (.A_N(_0339_),
    .B(_0345_),
    .Y(_0346_));
 sky130_fd_sc_hd__a21oi_1 _1142_ (.A1(_0317_),
    .A2(\MAC.add.b1[12] ),
    .B1(_0339_),
    .Y(_0347_));
 sky130_fd_sc_hd__a21o_1 _1143_ (.A1(_0345_),
    .A2(_0347_),
    .B1(_0338_),
    .X(_0348_));
 sky130_fd_sc_hd__a211o_1 _1144_ (.A1(_0345_),
    .A2(_0347_),
    .B1(_0336_),
    .C1(_0338_),
    .X(_0349_));
 sky130_fd_sc_hd__a31o_1 _1145_ (.A1(_0333_),
    .A2(_0337_),
    .A3(_0349_),
    .B1(_0334_),
    .X(_0350_));
 sky130_fd_sc_hd__a31oi_1 _1146_ (.A1(_0333_),
    .A2(_0337_),
    .A3(_0349_),
    .B1(_0334_),
    .Y(_0351_));
 sky130_fd_sc_hd__mux2_1 _1147_ (.A0(\MAC.add.b1[5] ),
    .A1(\MAC.add.a1[5] ),
    .S(net29),
    .X(_0352_));
 sky130_fd_sc_hd__xor2_2 _1148_ (.A(\MAC.add.a1[12] ),
    .B(\MAC.add.b1[12] ),
    .X(_0353_));
 sky130_fd_sc_hd__or2_1 _1149_ (.A(\MAC.add.a1[9] ),
    .B(_0318_),
    .X(_0354_));
 sky130_fd_sc_hd__xor2_2 _1150_ (.A(\MAC.add.a1[10] ),
    .B(\MAC.add.b1[10] ),
    .X(_0355_));
 sky130_fd_sc_hd__xnor2_2 _1151_ (.A(\MAC.add.a1[9] ),
    .B(\MAC.add.b1[9] ),
    .Y(_0356_));
 sky130_fd_sc_hd__xor2_2 _1152_ (.A(\MAC.add.a1[9] ),
    .B(\MAC.add.b1[9] ),
    .X(_0357_));
 sky130_fd_sc_hd__nor2_1 _1153_ (.A(_0355_),
    .B(_0357_),
    .Y(_0358_));
 sky130_fd_sc_hd__o31ai_2 _1154_ (.A1(_0341_),
    .A2(_0342_),
    .A3(_0356_),
    .B1(_0340_),
    .Y(_0359_));
 sky130_fd_sc_hd__o21ai_1 _1155_ (.A1(_0339_),
    .A2(_0359_),
    .B1(_0343_),
    .Y(_0360_));
 sky130_fd_sc_hd__or4_1 _1156_ (.A(\MAC.add.a1[10] ),
    .B(\MAC.add.a1[9] ),
    .C(\MAC.add.a1[14] ),
    .D(\MAC.add.a1[13] ),
    .X(_0361_));
 sky130_fd_sc_hd__nor3_1 _1157_ (.A(\MAC.add.a1[12] ),
    .B(\MAC.add.a1[11] ),
    .C(_0361_),
    .Y(_0362_));
 sky130_fd_sc_hd__or4_1 _1158_ (.A(\MAC.add.b1[10] ),
    .B(\MAC.add.b1[9] ),
    .C(\MAC.add.b1[14] ),
    .D(\MAC.add.b1[13] ),
    .X(_0363_));
 sky130_fd_sc_hd__nor3_1 _1159_ (.A(\MAC.add.b1[12] ),
    .B(\MAC.add.b1[11] ),
    .C(_0363_),
    .Y(_0364_));
 sky130_fd_sc_hd__nor2_1 _1160_ (.A(_0362_),
    .B(_0364_),
    .Y(_0365_));
 sky130_fd_sc_hd__or2_1 _1161_ (.A(_0362_),
    .B(_0364_),
    .X(_0366_));
 sky130_fd_sc_hd__xnor2_1 _1162_ (.A(_0353_),
    .B(_0360_),
    .Y(_0367_));
 sky130_fd_sc_hd__xnor2_1 _1163_ (.A(_0346_),
    .B(_0353_),
    .Y(_0368_));
 sky130_fd_sc_hd__mux2_1 _1164_ (.A0(_0367_),
    .A1(_0368_),
    .S(net28),
    .X(_0369_));
 sky130_fd_sc_hd__and2_1 _1165_ (.A(net32),
    .B(_0369_),
    .X(_0370_));
 sky130_fd_sc_hd__and2b_1 _1166_ (.A_N(_0336_),
    .B(_0337_),
    .X(_0371_));
 sky130_fd_sc_hd__nor4_1 _1167_ (.A(_0344_),
    .B(_0353_),
    .C(_0355_),
    .D(_0357_),
    .Y(_0372_));
 sky130_fd_sc_hd__or4_1 _1168_ (.A(_0344_),
    .B(_0353_),
    .C(_0355_),
    .D(_0357_),
    .X(_0373_));
 sky130_fd_sc_hd__a211o_1 _1169_ (.A1(_0345_),
    .A2(_0347_),
    .B1(_0372_),
    .C1(_0338_),
    .X(_0374_));
 sky130_fd_sc_hd__xor2_1 _1170_ (.A(_0371_),
    .B(_0374_),
    .X(_0375_));
 sky130_fd_sc_hd__a21oi_1 _1171_ (.A1(net28),
    .A2(_0373_),
    .B1(_0375_),
    .Y(_0376_));
 sky130_fd_sc_hd__a31o_1 _1172_ (.A1(net27),
    .A2(_0373_),
    .A3(_0375_),
    .B1(_0366_),
    .X(_0377_));
 sky130_fd_sc_hd__or2_1 _1173_ (.A(_0376_),
    .B(_0377_),
    .X(_0378_));
 sky130_fd_sc_hd__xnor2_1 _1174_ (.A(_0344_),
    .B(_0359_),
    .Y(_0379_));
 sky130_fd_sc_hd__o21ai_1 _1175_ (.A1(_0350_),
    .A2(_0358_),
    .B1(_0379_),
    .Y(_0380_));
 sky130_fd_sc_hd__o31a_1 _1176_ (.A1(net29),
    .A2(_0358_),
    .A3(_0379_),
    .B1(net32),
    .X(_0381_));
 sky130_fd_sc_hd__and2_2 _1177_ (.A(_0380_),
    .B(_0381_),
    .X(_0382_));
 sky130_fd_sc_hd__nand2_2 _1178_ (.A(_0380_),
    .B(_0381_),
    .Y(_0383_));
 sky130_fd_sc_hd__o2bb2a_2 _1179_ (.A1_N(net32),
    .A2_N(_0369_),
    .B1(_0376_),
    .B2(_0377_),
    .X(_0384_));
 sky130_fd_sc_hd__nand2b_1 _1180_ (.A_N(_0370_),
    .B(_0378_),
    .Y(_0385_));
 sky130_fd_sc_hd__nand2_1 _1181_ (.A(_0383_),
    .B(_0384_),
    .Y(_0386_));
 sky130_fd_sc_hd__xnor2_1 _1182_ (.A(_0354_),
    .B(_0355_),
    .Y(_0387_));
 sky130_fd_sc_hd__a311o_1 _1183_ (.A1(_0333_),
    .A2(_0337_),
    .A3(_0349_),
    .B1(_0356_),
    .C1(_0334_),
    .X(_0388_));
 sky130_fd_sc_hd__xnor2_1 _1184_ (.A(_0387_),
    .B(_0388_),
    .Y(_0389_));
 sky130_fd_sc_hd__and2_1 _1185_ (.A(net32),
    .B(_0389_),
    .X(_0390_));
 sky130_fd_sc_hd__nand2_1 _1186_ (.A(net32),
    .B(_0389_),
    .Y(_0391_));
 sky130_fd_sc_hd__o311ai_4 _1187_ (.A1(_0336_),
    .A2(_0348_),
    .A3(net33),
    .B1(_0337_),
    .C1(_0334_),
    .Y(_0392_));
 sky130_fd_sc_hd__a21o_1 _1188_ (.A1(_0337_),
    .A2(_0349_),
    .B1(_0333_),
    .X(_0393_));
 sky130_fd_sc_hd__or2_2 _1189_ (.A(\MAC.add.a1[14] ),
    .B(\MAC.add.b1[14] ),
    .X(_0394_));
 sky130_fd_sc_hd__a31oi_2 _1190_ (.A1(_0356_),
    .A2(_0392_),
    .A3(_0393_),
    .B1(_0366_),
    .Y(_0395_));
 sky130_fd_sc_hd__inv_2 _1191_ (.A(_0395_),
    .Y(_0396_));
 sky130_fd_sc_hd__or3_2 _1192_ (.A(_0386_),
    .B(_0390_),
    .C(_0395_),
    .X(_0397_));
 sky130_fd_sc_hd__inv_2 _1193_ (.A(_0397_),
    .Y(_0398_));
 sky130_fd_sc_hd__and3_1 _1194_ (.A(net32),
    .B(_0392_),
    .C(_0393_),
    .X(_0399_));
 sky130_fd_sc_hd__mux2_1 _1195_ (.A0(\MAC.add.b1[8] ),
    .A1(\MAC.add.a1[8] ),
    .S(net27),
    .X(_0400_));
 sky130_fd_sc_hd__o21a_1 _1196_ (.A1(_0357_),
    .A2(_0400_),
    .B1(_0399_),
    .X(_0401_));
 sky130_fd_sc_hd__nand2_1 _1197_ (.A(net26),
    .B(_0401_),
    .Y(_0402_));
 sky130_fd_sc_hd__mux2_1 _1198_ (.A0(\MAC.add.b1[8] ),
    .A1(\MAC.add.a1[8] ),
    .S(net29),
    .X(_0403_));
 sky130_fd_sc_hd__and4_2 _1199_ (.A(_0356_),
    .B(net32),
    .C(_0392_),
    .D(_0393_),
    .X(_0404_));
 sky130_fd_sc_hd__mux2_1 _1200_ (.A0(\MAC.add.b1[7] ),
    .A1(\MAC.add.a1[7] ),
    .S(net27),
    .X(_0405_));
 sky130_fd_sc_hd__and4_2 _1201_ (.A(_0357_),
    .B(net32),
    .C(_0392_),
    .D(_0393_),
    .X(_0406_));
 sky130_fd_sc_hd__a22o_1 _1202_ (.A1(_0404_),
    .A2(_0405_),
    .B1(_0406_),
    .B2(_0400_),
    .X(_0407_));
 sky130_fd_sc_hd__and3_1 _1203_ (.A(net32),
    .B(_0389_),
    .C(_0395_),
    .X(_0408_));
 sky130_fd_sc_hd__o21bai_1 _1204_ (.A1(_0390_),
    .A2(_0407_),
    .B1_N(_0408_),
    .Y(_0409_));
 sky130_fd_sc_hd__or2_1 _1205_ (.A(_0386_),
    .B(_0409_),
    .X(_0410_));
 sky130_fd_sc_hd__inv_2 _1206_ (.A(_0410_),
    .Y(_0411_));
 sky130_fd_sc_hd__mux2_1 _1207_ (.A0(\MAC.add.b1[7] ),
    .A1(\MAC.add.a1[7] ),
    .S(_0350_),
    .X(_0412_));
 sky130_fd_sc_hd__mux2_1 _1208_ (.A0(\MAC.add.b1[6] ),
    .A1(\MAC.add.a1[6] ),
    .S(net27),
    .X(_0413_));
 sky130_fd_sc_hd__a22o_1 _1209_ (.A1(_0405_),
    .A2(_0406_),
    .B1(_0413_),
    .B2(_0404_),
    .X(_0414_));
 sky130_fd_sc_hd__mux2_1 _1210_ (.A0(_0401_),
    .A1(_0414_),
    .S(net26),
    .X(_0415_));
 sky130_fd_sc_hd__nand2b_1 _1211_ (.A_N(_0386_),
    .B(_0415_),
    .Y(_0416_));
 sky130_fd_sc_hd__inv_2 _1212_ (.A(_0416_),
    .Y(_0417_));
 sky130_fd_sc_hd__mux2_1 _1213_ (.A0(\MAC.add.b1[6] ),
    .A1(\MAC.add.a1[6] ),
    .S(net29),
    .X(_0418_));
 sky130_fd_sc_hd__o22a_1 _1214_ (.A1(_0410_),
    .A2(_0412_),
    .B1(_0416_),
    .B2(_0418_),
    .X(_0419_));
 sky130_fd_sc_hd__mux2_1 _1215_ (.A0(\MAC.add.b1[5] ),
    .A1(\MAC.add.a1[5] ),
    .S(net27),
    .X(_0420_));
 sky130_fd_sc_hd__a22o_1 _1216_ (.A1(_0406_),
    .A2(_0413_),
    .B1(_0420_),
    .B2(_0404_),
    .X(_0421_));
 sky130_fd_sc_hd__mux2_1 _1217_ (.A0(_0407_),
    .A1(_0421_),
    .S(net26),
    .X(_0422_));
 sky130_fd_sc_hd__a21o_1 _1218_ (.A1(net26),
    .A2(_0396_),
    .B1(_0383_),
    .X(_0423_));
 sky130_fd_sc_hd__o211ai_2 _1219_ (.A1(_0382_),
    .A2(_0422_),
    .B1(_0423_),
    .C1(_0384_),
    .Y(_0424_));
 sky130_fd_sc_hd__inv_2 _1220_ (.A(_0424_),
    .Y(_0425_));
 sky130_fd_sc_hd__a22o_1 _1221_ (.A1(_0416_),
    .A2(_0418_),
    .B1(_0424_),
    .B2(_0352_),
    .X(_0426_));
 sky130_fd_sc_hd__mux2_1 _1222_ (.A0(\MAC.add.b1[4] ),
    .A1(\MAC.add.a1[4] ),
    .S(net27),
    .X(_0427_));
 sky130_fd_sc_hd__a22o_1 _1223_ (.A1(_0406_),
    .A2(_0420_),
    .B1(_0427_),
    .B2(_0404_),
    .X(_0428_));
 sky130_fd_sc_hd__mux2_1 _1224_ (.A0(_0414_),
    .A1(_0428_),
    .S(net26),
    .X(_0429_));
 sky130_fd_sc_hd__a21o_1 _1225_ (.A1(net26),
    .A2(_0401_),
    .B1(_0383_),
    .X(_0430_));
 sky130_fd_sc_hd__o211a_1 _1226_ (.A1(_0382_),
    .A2(_0429_),
    .B1(_0430_),
    .C1(_0384_),
    .X(_0431_));
 sky130_fd_sc_hd__mux2_1 _1227_ (.A0(\MAC.add.b1[4] ),
    .A1(\MAC.add.a1[4] ),
    .S(net29),
    .X(_0432_));
 sky130_fd_sc_hd__inv_2 _1228_ (.A(_0432_),
    .Y(_0433_));
 sky130_fd_sc_hd__a2bb2o_1 _1229_ (.A1_N(_0352_),
    .A2_N(_0424_),
    .B1(_0431_),
    .B2(_0433_),
    .X(_0434_));
 sky130_fd_sc_hd__a41o_1 _1230_ (.A1(_0378_),
    .A2(_0383_),
    .A3(net26),
    .A4(_0396_),
    .B1(_0384_),
    .X(_0435_));
 sky130_fd_sc_hd__mux2_1 _1231_ (.A0(\MAC.add.b1[3] ),
    .A1(\MAC.add.a1[3] ),
    .S(net27),
    .X(_0436_));
 sky130_fd_sc_hd__a22o_1 _1232_ (.A1(_0406_),
    .A2(_0427_),
    .B1(_0436_),
    .B2(_0404_),
    .X(_0437_));
 sky130_fd_sc_hd__or2_1 _1233_ (.A(net26),
    .B(_0437_),
    .X(_0438_));
 sky130_fd_sc_hd__mux2_1 _1234_ (.A0(\MAC.add.b1[1] ),
    .A1(\MAC.add.a1[1] ),
    .S(net27),
    .X(_0439_));
 sky130_fd_sc_hd__and2_1 _1235_ (.A(_0404_),
    .B(_0439_),
    .X(_0440_));
 sky130_fd_sc_hd__mux2_1 _1236_ (.A0(\MAC.add.b1[2] ),
    .A1(\MAC.add.a1[2] ),
    .S(net27),
    .X(_0441_));
 sky130_fd_sc_hd__and2_1 _1237_ (.A(_0406_),
    .B(_0441_),
    .X(_0442_));
 sky130_fd_sc_hd__o31a_1 _1238_ (.A1(_0390_),
    .A2(_0440_),
    .A3(_0442_),
    .B1(_0383_),
    .X(_0443_));
 sky130_fd_sc_hd__a221o_1 _1239_ (.A1(_0382_),
    .A2(_0422_),
    .B1(_0438_),
    .B2(_0443_),
    .C1(_0370_),
    .X(_0444_));
 sky130_fd_sc_hd__and2_1 _1240_ (.A(_0435_),
    .B(_0444_),
    .X(_0445_));
 sky130_fd_sc_hd__mux2_1 _1241_ (.A0(\MAC.add.b1[1] ),
    .A1(\MAC.add.a1[1] ),
    .S(net29),
    .X(_0446_));
 sky130_fd_sc_hd__inv_2 _1242_ (.A(_0446_),
    .Y(_0447_));
 sky130_fd_sc_hd__mux2_1 _1243_ (.A0(\MAC.add.b1[0] ),
    .A1(\MAC.add.a1[0] ),
    .S(net29),
    .X(_0448_));
 sky130_fd_sc_hd__mux2_1 _1244_ (.A0(\MAC.add.b1[0] ),
    .A1(\MAC.add.a1[0] ),
    .S(net27),
    .X(_0449_));
 sky130_fd_sc_hd__a22o_1 _1245_ (.A1(_0406_),
    .A2(_0439_),
    .B1(_0449_),
    .B2(_0404_),
    .X(_0450_));
 sky130_fd_sc_hd__or2_1 _1246_ (.A(_0370_),
    .B(_0382_),
    .X(_0451_));
 sky130_fd_sc_hd__a22o_1 _1247_ (.A1(_0406_),
    .A2(_0436_),
    .B1(_0441_),
    .B2(_0404_),
    .X(_0452_));
 sky130_fd_sc_hd__mux2_1 _1248_ (.A0(_0450_),
    .A1(_0452_),
    .S(_0390_),
    .X(_0453_));
 sky130_fd_sc_hd__a41o_1 _1249_ (.A1(_0378_),
    .A2(_0383_),
    .A3(net26),
    .A4(_0401_),
    .B1(_0384_),
    .X(_0454_));
 sky130_fd_sc_hd__o221a_1 _1250_ (.A1(_0383_),
    .A2(_0429_),
    .B1(_0451_),
    .B2(_0453_),
    .C1(_0454_),
    .X(_0455_));
 sky130_fd_sc_hd__a31oi_1 _1251_ (.A1(_0435_),
    .A2(_0444_),
    .A3(_0447_),
    .B1(_0455_),
    .Y(_0456_));
 sky130_fd_sc_hd__a21oi_1 _1252_ (.A1(_0435_),
    .A2(_0444_),
    .B1(_0447_),
    .Y(_0457_));
 sky130_fd_sc_hd__and2_1 _1253_ (.A(net26),
    .B(_0452_),
    .X(_0458_));
 sky130_fd_sc_hd__a21o_1 _1254_ (.A1(_0390_),
    .A2(_0428_),
    .B1(_0382_),
    .X(_0459_));
 sky130_fd_sc_hd__o221a_1 _1255_ (.A1(_0383_),
    .A2(_0415_),
    .B1(_0458_),
    .B2(_0459_),
    .C1(_0384_),
    .X(_0460_));
 sky130_fd_sc_hd__inv_2 _1256_ (.A(_0460_),
    .Y(_0461_));
 sky130_fd_sc_hd__mux2_1 _1257_ (.A0(\MAC.add.b1[2] ),
    .A1(\MAC.add.a1[2] ),
    .S(net29),
    .X(_0462_));
 sky130_fd_sc_hd__a221o_1 _1258_ (.A1(_0448_),
    .A2(_0456_),
    .B1(_0461_),
    .B2(_0462_),
    .C1(_0457_),
    .X(_0463_));
 sky130_fd_sc_hd__mux2_1 _1259_ (.A0(_0421_),
    .A1(_0437_),
    .S(_0391_),
    .X(_0464_));
 sky130_fd_sc_hd__nor2_1 _1260_ (.A(_0382_),
    .B(_0464_),
    .Y(_0465_));
 sky130_fd_sc_hd__a211oi_1 _1261_ (.A1(_0382_),
    .A2(_0409_),
    .B1(_0465_),
    .C1(_0385_),
    .Y(_0466_));
 sky130_fd_sc_hd__a211o_1 _1262_ (.A1(_0382_),
    .A2(_0409_),
    .B1(_0465_),
    .C1(_0385_),
    .X(_0467_));
 sky130_fd_sc_hd__mux2_1 _1263_ (.A0(\MAC.add.b1[3] ),
    .A1(\MAC.add.a1[3] ),
    .S(net29),
    .X(_0468_));
 sky130_fd_sc_hd__o22a_1 _1264_ (.A1(_0461_),
    .A2(_0462_),
    .B1(_0467_),
    .B2(_0468_),
    .X(_0469_));
 sky130_fd_sc_hd__and2_1 _1265_ (.A(_0410_),
    .B(_0412_),
    .X(_0470_));
 sky130_fd_sc_hd__or3_1 _1266_ (.A(_0397_),
    .B(_0402_),
    .C(_0403_),
    .X(_0471_));
 sky130_fd_sc_hd__nand2b_1 _1267_ (.A_N(_0426_),
    .B(_0434_),
    .Y(_0472_));
 sky130_fd_sc_hd__a21o_1 _1268_ (.A1(_0419_),
    .A2(_0472_),
    .B1(_0470_),
    .X(_0473_));
 sky130_fd_sc_hd__o21ai_1 _1269_ (.A1(_0431_),
    .A2(_0433_),
    .B1(_0419_),
    .Y(_0474_));
 sky130_fd_sc_hd__a211o_1 _1270_ (.A1(_0467_),
    .A2(_0468_),
    .B1(_0426_),
    .C1(_0434_),
    .X(_0475_));
 sky130_fd_sc_hd__a2111o_1 _1271_ (.A1(_0463_),
    .A2(_0469_),
    .B1(_0470_),
    .C1(_0474_),
    .D1(_0475_),
    .X(_0476_));
 sky130_fd_sc_hd__a221o_1 _1272_ (.A1(_0402_),
    .A2(_0403_),
    .B1(_0473_),
    .B2(_0476_),
    .C1(_0397_),
    .X(_0477_));
 sky130_fd_sc_hd__and2_1 _1273_ (.A(_0471_),
    .B(_0477_),
    .X(_0478_));
 sky130_fd_sc_hd__mux2_1 _1274_ (.A0(_0352_),
    .A1(_0425_),
    .S(net22),
    .X(_0479_));
 sky130_fd_sc_hd__mux2_1 _1275_ (.A0(_0468_),
    .A1(_0466_),
    .S(net21),
    .X(_0480_));
 sky130_fd_sc_hd__mux2_2 _1276_ (.A0(_0462_),
    .A1(_0460_),
    .S(net21),
    .X(_0481_));
 sky130_fd_sc_hd__and3_1 _1277_ (.A(_0455_),
    .B(_0471_),
    .C(_0477_),
    .X(_0482_));
 sky130_fd_sc_hd__a21boi_1 _1278_ (.A1(_0471_),
    .A2(_0477_),
    .B1_N(_0448_),
    .Y(_0483_));
 sky130_fd_sc_hd__or2_1 _1279_ (.A(_0482_),
    .B(_0483_),
    .X(_0484_));
 sky130_fd_sc_hd__a21oi_1 _1280_ (.A1(_0471_),
    .A2(_0477_),
    .B1(_0447_),
    .Y(_0485_));
 sky130_fd_sc_hd__and3_1 _1281_ (.A(_0445_),
    .B(_0471_),
    .C(_0477_),
    .X(_0486_));
 sky130_fd_sc_hd__or2_1 _1282_ (.A(_0485_),
    .B(_0486_),
    .X(_0487_));
 sky130_fd_sc_hd__or4_2 _1283_ (.A(_0482_),
    .B(_0483_),
    .C(_0485_),
    .D(_0486_),
    .X(_0488_));
 sky130_fd_sc_hd__or3_1 _1284_ (.A(_0480_),
    .B(_0481_),
    .C(_0488_),
    .X(_0489_));
 sky130_fd_sc_hd__mux2_2 _1285_ (.A0(_0432_),
    .A1(_0431_),
    .S(net21),
    .X(_0490_));
 sky130_fd_sc_hd__or2_1 _1286_ (.A(_0479_),
    .B(_0490_),
    .X(_0491_));
 sky130_fd_sc_hd__mux2_1 _1287_ (.A0(_0418_),
    .A1(_0417_),
    .S(net21),
    .X(_0492_));
 sky130_fd_sc_hd__mux2_1 _1288_ (.A0(_0412_),
    .A1(_0411_),
    .S(net21),
    .X(_0493_));
 sky130_fd_sc_hd__or4_1 _1289_ (.A(_0489_),
    .B(_0491_),
    .C(_0492_),
    .D(_0493_),
    .X(_0494_));
 sky130_fd_sc_hd__nor2_1 _1290_ (.A(_0386_),
    .B(_0402_),
    .Y(_0495_));
 sky130_fd_sc_hd__o31a_1 _1291_ (.A1(_0398_),
    .A2(_0494_),
    .A3(_0495_),
    .B1(net34),
    .X(_0496_));
 sky130_fd_sc_hd__mux2_2 _1292_ (.A0(_0403_),
    .A1(_0495_),
    .S(net22),
    .X(_0497_));
 sky130_fd_sc_hd__and2_1 _1293_ (.A(_0332_),
    .B(_0494_),
    .X(_0498_));
 sky130_fd_sc_hd__xor2_4 _1294_ (.A(_0497_),
    .B(_0498_),
    .X(_0499_));
 sky130_fd_sc_hd__mux2_2 _1295_ (.A0(_0495_),
    .A1(_0403_),
    .S(net21),
    .X(_0500_));
 sky130_fd_sc_hd__nand2_1 _1296_ (.A(_0499_),
    .B(_0500_),
    .Y(_0501_));
 sky130_fd_sc_hd__xnor2_4 _1297_ (.A(_0499_),
    .B(_0500_),
    .Y(_0502_));
 sky130_fd_sc_hd__and2_1 _1298_ (.A(net34),
    .B(_0489_),
    .X(_0503_));
 sky130_fd_sc_hd__o41a_1 _1299_ (.A1(_0480_),
    .A2(_0481_),
    .A3(_0488_),
    .A4(_0490_),
    .B1(net34),
    .X(_0504_));
 sky130_fd_sc_hd__xnor2_1 _1300_ (.A(_0479_),
    .B(_0504_),
    .Y(_0505_));
 sky130_fd_sc_hd__mux2_1 _1301_ (.A0(_0425_),
    .A1(_0352_),
    .S(net22),
    .X(_0506_));
 sky130_fd_sc_hd__inv_2 _1302_ (.A(_0506_),
    .Y(_0507_));
 sky130_fd_sc_hd__or2_1 _1303_ (.A(_0505_),
    .B(_0507_),
    .X(_0508_));
 sky130_fd_sc_hd__and2_1 _1304_ (.A(_0505_),
    .B(_0507_),
    .X(_0509_));
 sky130_fd_sc_hd__nand2_1 _1305_ (.A(_0505_),
    .B(_0507_),
    .Y(_0510_));
 sky130_fd_sc_hd__nand2_2 _1306_ (.A(_0508_),
    .B(_0510_),
    .Y(_0511_));
 sky130_fd_sc_hd__xnor2_4 _1307_ (.A(_0490_),
    .B(_0503_),
    .Y(_0512_));
 sky130_fd_sc_hd__mux2_2 _1308_ (.A0(_0431_),
    .A1(_0432_),
    .S(net22),
    .X(_0513_));
 sky130_fd_sc_hd__nand2b_1 _1309_ (.A_N(_0512_),
    .B(_0513_),
    .Y(_0514_));
 sky130_fd_sc_hd__xor2_4 _1310_ (.A(_0512_),
    .B(_0513_),
    .X(_0515_));
 sky130_fd_sc_hd__o21a_1 _1311_ (.A1(_0481_),
    .A2(_0488_),
    .B1(net34),
    .X(_0516_));
 sky130_fd_sc_hd__xor2_1 _1312_ (.A(_0480_),
    .B(_0516_),
    .X(_0517_));
 sky130_fd_sc_hd__mux2_1 _1313_ (.A0(_0466_),
    .A1(_0468_),
    .S(net22),
    .X(_0518_));
 sky130_fd_sc_hd__and2_1 _1314_ (.A(_0517_),
    .B(_0518_),
    .X(_0519_));
 sky130_fd_sc_hd__nor2_1 _1315_ (.A(_0517_),
    .B(_0518_),
    .Y(_0520_));
 sky130_fd_sc_hd__nand2_1 _1316_ (.A(net34),
    .B(_0488_),
    .Y(_0521_));
 sky130_fd_sc_hd__xnor2_2 _1317_ (.A(_0481_),
    .B(_0521_),
    .Y(_0522_));
 sky130_fd_sc_hd__mux2_1 _1318_ (.A0(_0460_),
    .A1(_0462_),
    .S(net21),
    .X(_0523_));
 sky130_fd_sc_hd__and2_1 _1319_ (.A(_0522_),
    .B(_0523_),
    .X(_0524_));
 sky130_fd_sc_hd__nand3_1 _1320_ (.A(net34),
    .B(_0484_),
    .C(_0487_),
    .Y(_0525_));
 sky130_fd_sc_hd__a21o_1 _1321_ (.A1(net34),
    .A2(_0484_),
    .B1(_0487_),
    .X(_0526_));
 sky130_fd_sc_hd__mux2_1 _1322_ (.A0(_0445_),
    .A1(_0446_),
    .S(net21),
    .X(_0527_));
 sky130_fd_sc_hd__and3_1 _1323_ (.A(_0525_),
    .B(_0526_),
    .C(_0527_),
    .X(_0528_));
 sky130_fd_sc_hd__nand2_2 _1324_ (.A(_0448_),
    .B(_0455_),
    .Y(_0529_));
 sky130_fd_sc_hd__a21oi_1 _1325_ (.A1(_0525_),
    .A2(_0526_),
    .B1(_0527_),
    .Y(_0530_));
 sky130_fd_sc_hd__or2_2 _1326_ (.A(_0528_),
    .B(_0530_),
    .X(_0531_));
 sky130_fd_sc_hd__o21bai_2 _1327_ (.A1(_0529_),
    .A2(_0530_),
    .B1_N(_0528_),
    .Y(_0532_));
 sky130_fd_sc_hd__xor2_2 _1328_ (.A(_0522_),
    .B(_0523_),
    .X(_0533_));
 sky130_fd_sc_hd__a21oi_1 _1329_ (.A1(_0532_),
    .A2(_0533_),
    .B1(_0524_),
    .Y(_0534_));
 sky130_fd_sc_hd__a211oi_1 _1330_ (.A1(_0532_),
    .A2(_0533_),
    .B1(_0519_),
    .C1(_0524_),
    .Y(_0535_));
 sky130_fd_sc_hd__or2_1 _1331_ (.A(_0520_),
    .B(_0535_),
    .X(_0536_));
 sky130_fd_sc_hd__or4_2 _1332_ (.A(_0511_),
    .B(_0515_),
    .C(_0520_),
    .D(_0535_),
    .X(_0537_));
 sky130_fd_sc_hd__o31a_1 _1333_ (.A1(_0489_),
    .A2(_0491_),
    .A3(_0492_),
    .B1(net34),
    .X(_0538_));
 sky130_fd_sc_hd__xor2_1 _1334_ (.A(_0493_),
    .B(_0538_),
    .X(_0539_));
 sky130_fd_sc_hd__mux2_1 _1335_ (.A0(_0411_),
    .A1(_0412_),
    .S(net21),
    .X(_0540_));
 sky130_fd_sc_hd__nor2_1 _1336_ (.A(_0539_),
    .B(_0540_),
    .Y(_0541_));
 sky130_fd_sc_hd__o21a_1 _1337_ (.A1(_0489_),
    .A2(_0491_),
    .B1(net34),
    .X(_0542_));
 sky130_fd_sc_hd__xor2_1 _1338_ (.A(_0492_),
    .B(_0542_),
    .X(_0543_));
 sky130_fd_sc_hd__mux2_1 _1339_ (.A0(_0417_),
    .A1(_0418_),
    .S(net21),
    .X(_0544_));
 sky130_fd_sc_hd__nand2_2 _1340_ (.A(_0543_),
    .B(_0544_),
    .Y(_0545_));
 sky130_fd_sc_hd__and2_1 _1341_ (.A(_0539_),
    .B(_0540_),
    .X(_0546_));
 sky130_fd_sc_hd__o21a_1 _1342_ (.A1(_0509_),
    .A2(_0514_),
    .B1(_0508_),
    .X(_0547_));
 sky130_fd_sc_hd__o21ba_1 _1343_ (.A1(_0541_),
    .A2(_0545_),
    .B1_N(_0546_),
    .X(_0548_));
 sky130_fd_sc_hd__or2_1 _1344_ (.A(_0543_),
    .B(_0544_),
    .X(_0549_));
 sky130_fd_sc_hd__nand2_1 _1345_ (.A(_0545_),
    .B(_0549_),
    .Y(_0550_));
 sky130_fd_sc_hd__or2_1 _1346_ (.A(_0541_),
    .B(_0546_),
    .X(_0551_));
 sky130_fd_sc_hd__o21bai_1 _1347_ (.A1(_0546_),
    .A2(_0549_),
    .B1_N(_0541_),
    .Y(_0552_));
 sky130_fd_sc_hd__a31o_1 _1348_ (.A1(_0537_),
    .A2(_0547_),
    .A3(_0548_),
    .B1(_0552_),
    .X(_0553_));
 sky130_fd_sc_hd__a311o_1 _1349_ (.A1(_0537_),
    .A2(_0547_),
    .A3(_0548_),
    .B1(_0552_),
    .C1(_0502_),
    .X(_0554_));
 sky130_fd_sc_hd__o21ai_1 _1350_ (.A1(_0494_),
    .A2(_0497_),
    .B1(net34),
    .Y(_0555_));
 sky130_fd_sc_hd__xnor2_1 _1351_ (.A(_0397_),
    .B(_0555_),
    .Y(_0556_));
 sky130_fd_sc_hd__nand3_1 _1352_ (.A(_0501_),
    .B(_0554_),
    .C(_0556_),
    .Y(_0557_));
 sky130_fd_sc_hd__and3b_2 _1353_ (.A_N(_0496_),
    .B(_0557_),
    .C(_0365_),
    .X(_0558_));
 sky130_fd_sc_hd__or3b_4 _1354_ (.A(_0366_),
    .B(_0496_),
    .C_N(_0557_),
    .X(_0559_));
 sky130_fd_sc_hd__xor2_4 _1355_ (.A(_0529_),
    .B(_0531_),
    .X(_0560_));
 sky130_fd_sc_hd__inv_2 _1356_ (.A(_0560_),
    .Y(_0561_));
 sky130_fd_sc_hd__a21o_1 _1357_ (.A1(_0501_),
    .A2(_0554_),
    .B1(_0556_),
    .X(_0562_));
 sky130_fd_sc_hd__and3_1 _1358_ (.A(_0365_),
    .B(_0557_),
    .C(_0562_),
    .X(_0563_));
 sky130_fd_sc_hd__nand3_2 _1359_ (.A(net32),
    .B(_0557_),
    .C(_0562_),
    .Y(_0564_));
 sky130_fd_sc_hd__a21o_2 _1360_ (.A1(_0537_),
    .A2(_0547_),
    .B1(_0550_),
    .X(_0565_));
 sky130_fd_sc_hd__and3_1 _1361_ (.A(_0545_),
    .B(_0551_),
    .C(_0565_),
    .X(_0566_));
 sky130_fd_sc_hd__nand3_2 _1362_ (.A(_0545_),
    .B(_0551_),
    .C(_0565_),
    .Y(_0567_));
 sky130_fd_sc_hd__a21oi_1 _1363_ (.A1(_0545_),
    .A2(_0565_),
    .B1(_0551_),
    .Y(_0568_));
 sky130_fd_sc_hd__a21o_1 _1364_ (.A1(_0545_),
    .A2(_0565_),
    .B1(_0551_),
    .X(_0569_));
 sky130_fd_sc_hd__nand2_2 _1365_ (.A(_0567_),
    .B(_0569_),
    .Y(_0570_));
 sky130_fd_sc_hd__nand3_2 _1366_ (.A(_0537_),
    .B(_0547_),
    .C(_0550_),
    .Y(_0571_));
 sky130_fd_sc_hd__and2_1 _1367_ (.A(_0565_),
    .B(_0571_),
    .X(_0572_));
 sky130_fd_sc_hd__nand2_2 _1368_ (.A(_0565_),
    .B(_0571_),
    .Y(_0573_));
 sky130_fd_sc_hd__xor2_4 _1369_ (.A(_0502_),
    .B(_0553_),
    .X(_0574_));
 sky130_fd_sc_hd__nor2_1 _1370_ (.A(_0572_),
    .B(_0574_),
    .Y(_0575_));
 sky130_fd_sc_hd__o31a_2 _1371_ (.A1(_0515_),
    .A2(_0520_),
    .A3(_0535_),
    .B1(_0514_),
    .X(_0576_));
 sky130_fd_sc_hd__xor2_2 _1372_ (.A(_0511_),
    .B(_0576_),
    .X(_0577_));
 sky130_fd_sc_hd__xnor2_2 _1373_ (.A(_0511_),
    .B(_0576_),
    .Y(_0578_));
 sky130_fd_sc_hd__xor2_1 _1374_ (.A(_0515_),
    .B(_0536_),
    .X(_0579_));
 sky130_fd_sc_hd__xnor2_2 _1375_ (.A(_0515_),
    .B(_0536_),
    .Y(_0580_));
 sky130_fd_sc_hd__nor2_1 _1376_ (.A(_0519_),
    .B(_0520_),
    .Y(_0581_));
 sky130_fd_sc_hd__xnor2_2 _1377_ (.A(_0534_),
    .B(_0581_),
    .Y(_0582_));
 sky130_fd_sc_hd__inv_2 _1378_ (.A(_0582_),
    .Y(_0583_));
 sky130_fd_sc_hd__xor2_2 _1379_ (.A(_0532_),
    .B(_0533_),
    .X(_0584_));
 sky130_fd_sc_hd__inv_2 _1380_ (.A(_0584_),
    .Y(_0585_));
 sky130_fd_sc_hd__or2_1 _1381_ (.A(_0582_),
    .B(_0584_),
    .X(_0586_));
 sky130_fd_sc_hd__or2_1 _1382_ (.A(_0579_),
    .B(_0586_),
    .X(_0587_));
 sky130_fd_sc_hd__o2111a_2 _1383_ (.A1(_0577_),
    .A2(_0587_),
    .B1(_0563_),
    .C1(_0570_),
    .D1(_0575_),
    .X(_0588_));
 sky130_fd_sc_hd__inv_2 _1384_ (.A(_0588_),
    .Y(_0589_));
 sky130_fd_sc_hd__or2_1 _1385_ (.A(_0448_),
    .B(_0455_),
    .X(_0590_));
 sky130_fd_sc_hd__nand2_2 _1386_ (.A(_0529_),
    .B(_0590_),
    .Y(_0591_));
 sky130_fd_sc_hd__or2_1 _1387_ (.A(_0560_),
    .B(_0591_),
    .X(_0592_));
 sky130_fd_sc_hd__a21o_1 _1388_ (.A1(_0585_),
    .A2(_0592_),
    .B1(_0582_),
    .X(_0593_));
 sky130_fd_sc_hd__a21oi_1 _1389_ (.A1(_0580_),
    .A2(_0593_),
    .B1(_0577_),
    .Y(_0594_));
 sky130_fd_sc_hd__or3_1 _1390_ (.A(_0572_),
    .B(_0574_),
    .C(_0594_),
    .X(_0595_));
 sky130_fd_sc_hd__nand2_1 _1391_ (.A(_0563_),
    .B(_0595_),
    .Y(_0596_));
 sky130_fd_sc_hd__or3_1 _1392_ (.A(_0566_),
    .B(_0568_),
    .C(_0574_),
    .X(_0597_));
 sky130_fd_sc_hd__and3_2 _1393_ (.A(_0563_),
    .B(_0595_),
    .C(_0597_),
    .X(_0598_));
 sky130_fd_sc_hd__nor2_1 _1394_ (.A(_0591_),
    .B(_0598_),
    .Y(_0599_));
 sky130_fd_sc_hd__or3b_1 _1395_ (.A(_0577_),
    .B(_0579_),
    .C_N(_0586_),
    .X(_0600_));
 sky130_fd_sc_hd__a311oi_4 _1396_ (.A1(_0570_),
    .A2(_0573_),
    .A3(_0600_),
    .B1(_0574_),
    .C1(_0564_),
    .Y(_0601_));
 sky130_fd_sc_hd__or3_1 _1397_ (.A(_0591_),
    .B(_0598_),
    .C(net20),
    .X(_0602_));
 sky130_fd_sc_hd__a21o_1 _1398_ (.A1(_0567_),
    .A2(_0569_),
    .B1(_0574_),
    .X(_0603_));
 sky130_fd_sc_hd__a21oi_1 _1399_ (.A1(_0565_),
    .A2(_0571_),
    .B1(_0577_),
    .Y(_0604_));
 sky130_fd_sc_hd__nand2_1 _1400_ (.A(_0573_),
    .B(_0578_),
    .Y(_0605_));
 sky130_fd_sc_hd__a2111o_1 _1401_ (.A1(_0565_),
    .A2(_0571_),
    .B1(_0577_),
    .C1(_0579_),
    .D1(_0586_),
    .X(_0606_));
 sky130_fd_sc_hd__a211o_1 _1402_ (.A1(_0567_),
    .A2(_0569_),
    .B1(_0574_),
    .C1(_0606_),
    .X(_0607_));
 sky130_fd_sc_hd__nand2_1 _1403_ (.A(_0561_),
    .B(_0591_),
    .Y(_0608_));
 sky130_fd_sc_hd__nor3b_1 _1404_ (.A(_0564_),
    .B(_0607_),
    .C_N(_0608_),
    .Y(_0609_));
 sky130_fd_sc_hd__or2_2 _1405_ (.A(_0558_),
    .B(_0609_),
    .X(_0610_));
 sky130_fd_sc_hd__nor2_1 _1406_ (.A(_0602_),
    .B(_0610_),
    .Y(_0611_));
 sky130_fd_sc_hd__nor2_1 _1407_ (.A(_0588_),
    .B(_0609_),
    .Y(_0612_));
 sky130_fd_sc_hd__nor2_1 _1408_ (.A(_0588_),
    .B(_0610_),
    .Y(_0613_));
 sky130_fd_sc_hd__a22o_1 _1409_ (.A1(_0558_),
    .A2(_0560_),
    .B1(_0589_),
    .B2(_0611_),
    .X(_0614_));
 sky130_fd_sc_hd__mux2_1 _1410_ (.A0(\MAC.add.a1[9] ),
    .A1(\MAC.add.b1[9] ),
    .S(net28),
    .X(_0615_));
 sky130_fd_sc_hd__mux2_1 _1411_ (.A0(\MAC.add.a1[11] ),
    .A1(\MAC.add.b1[11] ),
    .S(net28),
    .X(_0616_));
 sky130_fd_sc_hd__mux2_1 _1412_ (.A0(\MAC.add.a1[10] ),
    .A1(\MAC.add.b1[10] ),
    .S(net28),
    .X(_0617_));
 sky130_fd_sc_hd__or3_1 _1413_ (.A(_0615_),
    .B(_0616_),
    .C(_0617_),
    .X(_0618_));
 sky130_fd_sc_hd__and4_2 _1414_ (.A(_0365_),
    .B(_0496_),
    .C(_0557_),
    .D(_0562_),
    .X(_0619_));
 sky130_fd_sc_hd__nor2_1 _1415_ (.A(_0587_),
    .B(_0592_),
    .Y(_0620_));
 sky130_fd_sc_hd__o31a_1 _1416_ (.A1(_0603_),
    .A2(_0605_),
    .A3(_0620_),
    .B1(_0619_),
    .X(_0621_));
 sky130_fd_sc_hd__or2_1 _1417_ (.A(_0616_),
    .B(_0621_),
    .X(_0622_));
 sky130_fd_sc_hd__o311a_1 _1418_ (.A1(_0603_),
    .A2(_0605_),
    .A3(_0620_),
    .B1(_0619_),
    .C1(_0616_),
    .X(_0623_));
 sky130_fd_sc_hd__nand2_1 _1419_ (.A(_0616_),
    .B(_0621_),
    .Y(_0624_));
 sky130_fd_sc_hd__o211ai_1 _1420_ (.A1(_0584_),
    .A2(_0592_),
    .B1(_0580_),
    .C1(_0583_),
    .Y(_0625_));
 sky130_fd_sc_hd__a221o_1 _1421_ (.A1(_0567_),
    .A2(_0569_),
    .B1(_0604_),
    .B2(_0625_),
    .C1(_0574_),
    .X(_0626_));
 sky130_fd_sc_hd__a21oi_1 _1422_ (.A1(_0619_),
    .A2(_0626_),
    .B1(_0617_),
    .Y(_0627_));
 sky130_fd_sc_hd__a21o_1 _1423_ (.A1(_0619_),
    .A2(_0626_),
    .B1(_0617_),
    .X(_0628_));
 sky130_fd_sc_hd__and3_1 _1424_ (.A(_0617_),
    .B(_0619_),
    .C(_0626_),
    .X(_0629_));
 sky130_fd_sc_hd__a31o_1 _1425_ (.A1(_0563_),
    .A2(_0595_),
    .A3(_0597_),
    .B1(_0558_),
    .X(_0630_));
 sky130_fd_sc_hd__nand2_1 _1426_ (.A(_0615_),
    .B(_0630_),
    .Y(_0631_));
 sky130_fd_sc_hd__nor2_1 _1427_ (.A(_0627_),
    .B(_0631_),
    .Y(_0632_));
 sky130_fd_sc_hd__a311o_1 _1428_ (.A1(_0615_),
    .A2(_0628_),
    .A3(_0630_),
    .B1(_0629_),
    .C1(_0623_),
    .X(_0633_));
 sky130_fd_sc_hd__nand2_1 _1429_ (.A(_0622_),
    .B(_0624_),
    .Y(_0634_));
 sky130_fd_sc_hd__nand2_1 _1430_ (.A(_0622_),
    .B(_0633_),
    .Y(_0635_));
 sky130_fd_sc_hd__a21bo_1 _1431_ (.A1(_0622_),
    .A2(_0633_),
    .B1_N(_0618_),
    .X(_0636_));
 sky130_fd_sc_hd__mux2_1 _1432_ (.A0(\MAC.add.a1[12] ),
    .A1(\MAC.add.b1[12] ),
    .S(net28),
    .X(_0637_));
 sky130_fd_sc_hd__or2_1 _1433_ (.A(_0618_),
    .B(_0637_),
    .X(_0638_));
 sky130_fd_sc_hd__nand2_1 _1434_ (.A(_0618_),
    .B(_0637_),
    .Y(_0639_));
 sky130_fd_sc_hd__nand2_1 _1435_ (.A(_0638_),
    .B(_0639_),
    .Y(_0640_));
 sky130_fd_sc_hd__o21a_1 _1436_ (.A1(_0560_),
    .A2(_0607_),
    .B1(_0619_),
    .X(_0641_));
 sky130_fd_sc_hd__o21a_1 _1437_ (.A1(_0607_),
    .A2(_0608_),
    .B1(_0619_),
    .X(_0642_));
 sky130_fd_sc_hd__mux2_2 _1438_ (.A0(\MAC.add.a1[13] ),
    .A1(\MAC.add.b1[13] ),
    .S(net28),
    .X(_0643_));
 sky130_fd_sc_hd__nor2_1 _1439_ (.A(_0638_),
    .B(_0643_),
    .Y(_0644_));
 sky130_fd_sc_hd__and2_1 _1440_ (.A(_0638_),
    .B(_0643_),
    .X(_0645_));
 sky130_fd_sc_hd__nor2_1 _1441_ (.A(_0644_),
    .B(_0645_),
    .Y(_0646_));
 sky130_fd_sc_hd__nor2_1 _1442_ (.A(_0642_),
    .B(_0646_),
    .Y(_0647_));
 sky130_fd_sc_hd__xnor2_1 _1443_ (.A(_0394_),
    .B(_0644_),
    .Y(_0648_));
 sky130_fd_sc_hd__o22a_1 _1444_ (.A1(_0640_),
    .A2(_0641_),
    .B1(_0647_),
    .B2(_0648_),
    .X(_0649_));
 sky130_fd_sc_hd__nand2_1 _1445_ (.A(_0642_),
    .B(_0646_),
    .Y(_0650_));
 sky130_fd_sc_hd__a2111o_1 _1446_ (.A1(_0648_),
    .A2(_0650_),
    .B1(_0394_),
    .C1(_0640_),
    .D1(_0643_),
    .X(_0651_));
 sky130_fd_sc_hd__a21oi_2 _1447_ (.A1(_0636_),
    .A2(_0649_),
    .B1(_0651_),
    .Y(_0652_));
 sky130_fd_sc_hd__and4_1 _1448_ (.A(\MAC.add.a1[14] ),
    .B(\MAC.add.a1[13] ),
    .C(\MAC.add.a1[15] ),
    .D(\MAC.add.a1[0] ),
    .X(_0653_));
 sky130_fd_sc_hd__and4_1 _1449_ (.A(\MAC.add.a1[12] ),
    .B(\MAC.add.a1[11] ),
    .C(\MAC.add.a1[10] ),
    .D(\MAC.add.a1[9] ),
    .X(_0654_));
 sky130_fd_sc_hd__and4_1 _1450_ (.A(\MAC.add.a1[5] ),
    .B(\MAC.add.a1[6] ),
    .C(\MAC.add.a1[7] ),
    .D(\MAC.add.a1[8] ),
    .X(_0655_));
 sky130_fd_sc_hd__and4_1 _1451_ (.A(\MAC.add.a1[1] ),
    .B(\MAC.add.a1[2] ),
    .C(\MAC.add.a1[3] ),
    .D(\MAC.add.a1[4] ),
    .X(_0656_));
 sky130_fd_sc_hd__and4_2 _1452_ (.A(_0653_),
    .B(_0654_),
    .C(_0655_),
    .D(_0656_),
    .X(_0657_));
 sky130_fd_sc_hd__and4_1 _1453_ (.A(\MAC.add.b1[14] ),
    .B(\MAC.add.b1[13] ),
    .C(\MAC.add.b1[15] ),
    .D(\MAC.add.b1[0] ),
    .X(_0658_));
 sky130_fd_sc_hd__and3_1 _1454_ (.A(\MAC.add.b1[12] ),
    .B(\MAC.add.b1[11] ),
    .C(\MAC.add.b1[10] ),
    .X(_0659_));
 sky130_fd_sc_hd__and3_1 _1455_ (.A(\MAC.add.b1[9] ),
    .B(_0658_),
    .C(_0659_),
    .X(_0660_));
 sky130_fd_sc_hd__and4_1 _1456_ (.A(\MAC.add.b1[1] ),
    .B(\MAC.add.b1[2] ),
    .C(\MAC.add.b1[3] ),
    .D(\MAC.add.b1[4] ),
    .X(_0661_));
 sky130_fd_sc_hd__and4_1 _1457_ (.A(\MAC.add.b1[5] ),
    .B(\MAC.add.b1[6] ),
    .C(\MAC.add.b1[7] ),
    .D(\MAC.add.b1[8] ),
    .X(_0662_));
 sky130_fd_sc_hd__a31o_1 _1458_ (.A1(_0660_),
    .A2(_0661_),
    .A3(_0662_),
    .B1(_0657_),
    .X(_0663_));
 sky130_fd_sc_hd__a31oi_4 _1459_ (.A1(_0660_),
    .A2(_0661_),
    .A3(_0662_),
    .B1(_0657_),
    .Y(_0664_));
 sky130_fd_sc_hd__a31o_1 _1460_ (.A1(_0660_),
    .A2(_0661_),
    .A3(_0662_),
    .B1(_0657_),
    .X(_0665_));
 sky130_fd_sc_hd__and4_1 _1461_ (.A(_0615_),
    .B(_0617_),
    .C(_0637_),
    .D(_0643_),
    .X(_0666_));
 sky130_fd_sc_hd__nand3_1 _1462_ (.A(_0394_),
    .B(_0616_),
    .C(_0666_),
    .Y(_0667_));
 sky130_fd_sc_hd__or2_4 _1463_ (.A(_0559_),
    .B(_0667_),
    .X(_0668_));
 sky130_fd_sc_hd__o31a_1 _1464_ (.A1(_0614_),
    .A2(net18),
    .A3(_0665_),
    .B1(_0668_),
    .X(\MAC.add.c_add[0] ));
 sky130_fd_sc_hd__mux2_1 _1465_ (.A0(_0561_),
    .A1(_0591_),
    .S(_0598_),
    .X(_0669_));
 sky130_fd_sc_hd__or2_1 _1466_ (.A(net20),
    .B(_0669_),
    .X(_0670_));
 sky130_fd_sc_hd__or3_1 _1467_ (.A(_0588_),
    .B(_0609_),
    .C(_0670_),
    .X(_0671_));
 sky130_fd_sc_hd__mux2_1 _1468_ (.A0(_0585_),
    .A1(_0671_),
    .S(_0559_),
    .X(_0672_));
 sky130_fd_sc_hd__o21ba_2 _1469_ (.A1(_0559_),
    .A2(_0667_),
    .B1_N(_0663_),
    .X(_0673_));
 sky130_fd_sc_hd__nand2_1 _1470_ (.A(_0672_),
    .B(_0673_),
    .Y(\MAC.add.c_add[1] ));
 sky130_fd_sc_hd__mux2_1 _1471_ (.A0(_0584_),
    .A1(_0560_),
    .S(_0598_),
    .X(_0674_));
 sky130_fd_sc_hd__mux2_1 _1472_ (.A0(_0674_),
    .A1(_0599_),
    .S(net20),
    .X(_0675_));
 sky130_fd_sc_hd__a22o_1 _1473_ (.A1(_0558_),
    .A2(_0582_),
    .B1(_0613_),
    .B2(_0675_),
    .X(_0676_));
 sky130_fd_sc_hd__nor2_1 _1474_ (.A(_0665_),
    .B(_0676_),
    .Y(_0677_));
 sky130_fd_sc_hd__o21ai_1 _1475_ (.A1(_0652_),
    .A2(_0677_),
    .B1(_0668_),
    .Y(\MAC.add.c_add[2] ));
 sky130_fd_sc_hd__mux2_1 _1476_ (.A0(_0583_),
    .A1(_0585_),
    .S(_0598_),
    .X(_0678_));
 sky130_fd_sc_hd__mux2_1 _1477_ (.A0(_0678_),
    .A1(_0669_),
    .S(_0601_),
    .X(_0679_));
 sky130_fd_sc_hd__or3_1 _1478_ (.A(_0588_),
    .B(_0610_),
    .C(_0679_),
    .X(_0680_));
 sky130_fd_sc_hd__o211a_1 _1479_ (.A1(_0559_),
    .A2(_0580_),
    .B1(_0664_),
    .C1(_0680_),
    .X(_0681_));
 sky130_fd_sc_hd__o21ai_1 _1480_ (.A1(net18),
    .A2(_0681_),
    .B1(_0668_),
    .Y(\MAC.add.c_add[3] ));
 sky130_fd_sc_hd__mux2_1 _1481_ (.A0(_0579_),
    .A1(_0582_),
    .S(_0598_),
    .X(_0682_));
 sky130_fd_sc_hd__mux2_1 _1482_ (.A0(_0682_),
    .A1(_0674_),
    .S(net20),
    .X(_0683_));
 sky130_fd_sc_hd__o22ai_1 _1483_ (.A1(_0611_),
    .A2(_0613_),
    .B1(_0683_),
    .B2(_0588_),
    .Y(_0684_));
 sky130_fd_sc_hd__o211a_1 _1484_ (.A1(_0559_),
    .A2(_0578_),
    .B1(_0664_),
    .C1(_0684_),
    .X(_0685_));
 sky130_fd_sc_hd__o21ai_1 _1485_ (.A1(net18),
    .A2(_0685_),
    .B1(_0668_),
    .Y(\MAC.add.c_add[4] ));
 sky130_fd_sc_hd__mux2_1 _1486_ (.A0(_0578_),
    .A1(_0580_),
    .S(_0598_),
    .X(_0686_));
 sky130_fd_sc_hd__mux2_1 _1487_ (.A0(_0686_),
    .A1(_0678_),
    .S(_0601_),
    .X(_0687_));
 sky130_fd_sc_hd__a211o_1 _1488_ (.A1(_0588_),
    .A2(_0670_),
    .B1(_0687_),
    .C1(_0610_),
    .X(_0688_));
 sky130_fd_sc_hd__o211a_1 _1489_ (.A1(_0559_),
    .A2(_0573_),
    .B1(_0664_),
    .C1(_0688_),
    .X(_0689_));
 sky130_fd_sc_hd__o21ai_1 _1490_ (.A1(net18),
    .A2(_0689_),
    .B1(_0668_),
    .Y(\MAC.add.c_add[5] ));
 sky130_fd_sc_hd__mux2_1 _1491_ (.A0(_0573_),
    .A1(_0578_),
    .S(_0598_),
    .X(_0690_));
 sky130_fd_sc_hd__nor2_1 _1492_ (.A(net20),
    .B(_0690_),
    .Y(_0691_));
 sky130_fd_sc_hd__a211o_1 _1493_ (.A1(net20),
    .A2(_0682_),
    .B1(_0691_),
    .C1(_0588_),
    .X(_0692_));
 sky130_fd_sc_hd__o21ba_1 _1494_ (.A1(_0589_),
    .A2(_0675_),
    .B1_N(_0610_),
    .X(_0693_));
 sky130_fd_sc_hd__o21ai_1 _1495_ (.A1(_0559_),
    .A2(_0570_),
    .B1(_0664_),
    .Y(_0694_));
 sky130_fd_sc_hd__a21oi_1 _1496_ (.A1(_0692_),
    .A2(_0693_),
    .B1(_0694_),
    .Y(_0695_));
 sky130_fd_sc_hd__o21ai_1 _1497_ (.A1(_0652_),
    .A2(_0695_),
    .B1(_0668_),
    .Y(\MAC.add.c_add[6] ));
 sky130_fd_sc_hd__a22o_1 _1498_ (.A1(_0570_),
    .A2(_0596_),
    .B1(_0598_),
    .B2(_0573_),
    .X(_0696_));
 sky130_fd_sc_hd__mux2_1 _1499_ (.A0(_0696_),
    .A1(_0686_),
    .S(_0601_),
    .X(_0697_));
 sky130_fd_sc_hd__o21a_1 _1500_ (.A1(_0589_),
    .A2(_0679_),
    .B1(_0559_),
    .X(_0698_));
 sky130_fd_sc_hd__a2bb2o_1 _1501_ (.A1_N(_0559_),
    .A2_N(_0574_),
    .B1(_0697_),
    .B2(_0698_),
    .X(_0699_));
 sky130_fd_sc_hd__a21oi_1 _1502_ (.A1(_0673_),
    .A2(_0699_),
    .B1(net18),
    .Y(\MAC.add.c_add[7] ));
 sky130_fd_sc_hd__nor2_1 _1503_ (.A(_0589_),
    .B(_0683_),
    .Y(_0700_));
 sky130_fd_sc_hd__o21a_1 _1504_ (.A1(_0558_),
    .A2(_0602_),
    .B1(_0610_),
    .X(_0701_));
 sky130_fd_sc_hd__nand2b_1 _1505_ (.A_N(_0690_),
    .B(net20),
    .Y(_0702_));
 sky130_fd_sc_hd__a21bo_1 _1506_ (.A1(_0563_),
    .A2(_0570_),
    .B1_N(_0574_),
    .X(_0703_));
 sky130_fd_sc_hd__a31o_1 _1507_ (.A1(_0612_),
    .A2(_0702_),
    .A3(_0703_),
    .B1(_0701_),
    .X(_0704_));
 sky130_fd_sc_hd__nand2_1 _1508_ (.A(_0558_),
    .B(_0564_),
    .Y(_0705_));
 sky130_fd_sc_hd__o211a_1 _1509_ (.A1(_0700_),
    .A2(_0704_),
    .B1(_0705_),
    .C1(_0664_),
    .X(_0706_));
 sky130_fd_sc_hd__o21ai_1 _1510_ (.A1(_0652_),
    .A2(_0706_),
    .B1(_0668_),
    .Y(\MAC.add.c_add[8] ));
 sky130_fd_sc_hd__or2_1 _1511_ (.A(_0615_),
    .B(_0630_),
    .X(_0707_));
 sky130_fd_sc_hd__and2_1 _1512_ (.A(_0631_),
    .B(_0707_),
    .X(_0708_));
 sky130_fd_sc_hd__o31a_1 _1513_ (.A1(net18),
    .A2(_0665_),
    .A3(_0708_),
    .B1(_0668_),
    .X(\MAC.add.c_add[9] ));
 sky130_fd_sc_hd__nor2_1 _1514_ (.A(_0627_),
    .B(_0629_),
    .Y(_0709_));
 sky130_fd_sc_hd__xor2_1 _1515_ (.A(_0631_),
    .B(_0709_),
    .X(_0710_));
 sky130_fd_sc_hd__a21o_1 _1516_ (.A1(_0664_),
    .A2(_0710_),
    .B1(net18),
    .X(_0711_));
 sky130_fd_sc_hd__nand2_1 _1517_ (.A(_0668_),
    .B(_0711_),
    .Y(\MAC.add.c_add[10] ));
 sky130_fd_sc_hd__o21ai_1 _1518_ (.A1(_0629_),
    .A2(_0632_),
    .B1(_0634_),
    .Y(_0712_));
 sky130_fd_sc_hd__o31a_1 _1519_ (.A1(_0629_),
    .A2(_0632_),
    .A3(_0634_),
    .B1(_0673_),
    .X(_0713_));
 sky130_fd_sc_hd__a21oi_1 _1520_ (.A1(_0712_),
    .A2(_0713_),
    .B1(net18),
    .Y(\MAC.add.c_add[11] ));
 sky130_fd_sc_hd__and2_1 _1521_ (.A(_0637_),
    .B(_0641_),
    .X(_0714_));
 sky130_fd_sc_hd__or2_1 _1522_ (.A(_0637_),
    .B(_0641_),
    .X(_0715_));
 sky130_fd_sc_hd__nand2b_1 _1523_ (.A_N(_0714_),
    .B(_0715_),
    .Y(_0716_));
 sky130_fd_sc_hd__xnor2_1 _1524_ (.A(_0635_),
    .B(_0716_),
    .Y(_0717_));
 sky130_fd_sc_hd__a21oi_1 _1525_ (.A1(_0673_),
    .A2(_0717_),
    .B1(_0652_),
    .Y(\MAC.add.c_add[12] ));
 sky130_fd_sc_hd__a31o_1 _1526_ (.A1(_0622_),
    .A2(_0633_),
    .A3(_0715_),
    .B1(_0714_),
    .X(_0718_));
 sky130_fd_sc_hd__and2_1 _1527_ (.A(_0642_),
    .B(_0643_),
    .X(_0719_));
 sky130_fd_sc_hd__or2_1 _1528_ (.A(_0642_),
    .B(_0643_),
    .X(_0720_));
 sky130_fd_sc_hd__and2b_1 _1529_ (.A_N(_0719_),
    .B(_0720_),
    .X(_0721_));
 sky130_fd_sc_hd__xnor2_1 _1530_ (.A(_0718_),
    .B(_0721_),
    .Y(_0722_));
 sky130_fd_sc_hd__a21oi_1 _1531_ (.A1(_0673_),
    .A2(_0722_),
    .B1(net18),
    .Y(\MAC.add.c_add[13] ));
 sky130_fd_sc_hd__a21o_1 _1532_ (.A1(_0718_),
    .A2(_0720_),
    .B1(_0719_),
    .X(_0723_));
 sky130_fd_sc_hd__xnor2_1 _1533_ (.A(_0394_),
    .B(_0642_),
    .Y(_0724_));
 sky130_fd_sc_hd__nand2_1 _1534_ (.A(_0723_),
    .B(_0724_),
    .Y(_0725_));
 sky130_fd_sc_hd__or2_1 _1535_ (.A(_0723_),
    .B(_0724_),
    .X(_0726_));
 sky130_fd_sc_hd__a31oi_1 _1536_ (.A1(_0673_),
    .A2(_0725_),
    .A3(_0726_),
    .B1(net18),
    .Y(\MAC.add.c_add[14] ));
 sky130_fd_sc_hd__and4_1 _1537_ (.A(_0333_),
    .B(_0335_),
    .C(_0371_),
    .D(_0372_),
    .X(_0727_));
 sky130_fd_sc_hd__nor2_1 _1538_ (.A(\MAC.add.b1[8] ),
    .B(_0327_),
    .Y(_0728_));
 sky130_fd_sc_hd__a2bb2o_1 _1539_ (.A1_N(_0324_),
    .A2_N(\MAC.add.a1[6] ),
    .B1(\MAC.add.b1[7] ),
    .B2(_0325_),
    .X(_0729_));
 sky130_fd_sc_hd__nor2_1 _1540_ (.A(\MAC.add.b1[7] ),
    .B(_0325_),
    .Y(_0730_));
 sky130_fd_sc_hd__a211o_1 _1541_ (.A1(_0324_),
    .A2(\MAC.add.a1[6] ),
    .B1(_0729_),
    .C1(_0730_),
    .X(_0731_));
 sky130_fd_sc_hd__a221o_1 _1542_ (.A1(_0321_),
    .A2(\MAC.add.a1[4] ),
    .B1(_0322_),
    .B2(\MAC.add.a1[5] ),
    .C1(_0731_),
    .X(_0732_));
 sky130_fd_sc_hd__and2b_1 _1543_ (.A_N(\MAC.add.b1[3] ),
    .B(\MAC.add.a1[3] ),
    .X(_0733_));
 sky130_fd_sc_hd__nor2_1 _1544_ (.A(\MAC.add.a1[2] ),
    .B(_0733_),
    .Y(_0734_));
 sky130_fd_sc_hd__and2b_1 _1545_ (.A_N(\MAC.add.a1[3] ),
    .B(\MAC.add.b1[3] ),
    .X(_0735_));
 sky130_fd_sc_hd__nor2_1 _1546_ (.A(_0321_),
    .B(\MAC.add.a1[4] ),
    .Y(_0736_));
 sky130_fd_sc_hd__a211oi_1 _1547_ (.A1(\MAC.add.b1[2] ),
    .A2(_0734_),
    .B1(_0735_),
    .C1(_0736_),
    .Y(_0737_));
 sky130_fd_sc_hd__xor2_1 _1548_ (.A(\MAC.add.b1[2] ),
    .B(\MAC.add.a1[2] ),
    .X(_0738_));
 sky130_fd_sc_hd__or3_1 _1549_ (.A(_0733_),
    .B(_0735_),
    .C(_0738_),
    .X(_0739_));
 sky130_fd_sc_hd__or3b_1 _1550_ (.A(\MAC.add.a1[1] ),
    .B(_0739_),
    .C_N(\MAC.add.b1[1] ),
    .X(_0740_));
 sky130_fd_sc_hd__xor2_1 _1551_ (.A(\MAC.add.b1[1] ),
    .B(\MAC.add.a1[1] ),
    .X(_0741_));
 sky130_fd_sc_hd__a211o_1 _1552_ (.A1(_0319_),
    .A2(\MAC.add.a1[0] ),
    .B1(_0739_),
    .C1(_0741_),
    .X(_0742_));
 sky130_fd_sc_hd__o21ai_1 _1553_ (.A1(\MAC.add.b1[7] ),
    .A2(_0325_),
    .B1(_0729_),
    .Y(_0743_));
 sky130_fd_sc_hd__a31o_1 _1554_ (.A1(_0737_),
    .A2(_0740_),
    .A3(_0742_),
    .B1(_0732_),
    .X(_0744_));
 sky130_fd_sc_hd__o32a_1 _1555_ (.A1(_0322_),
    .A2(\MAC.add.a1[5] ),
    .A3(_0731_),
    .B1(\MAC.add.a1[8] ),
    .B2(_0326_),
    .X(_0745_));
 sky130_fd_sc_hd__a31o_1 _1556_ (.A1(_0743_),
    .A2(_0744_),
    .A3(_0745_),
    .B1(_0728_),
    .X(_0746_));
 sky130_fd_sc_hd__a221o_1 _1557_ (.A1(\MAC.add.b1[0] ),
    .A2(_0320_),
    .B1(\MAC.add.b1[8] ),
    .B2(_0327_),
    .C1(_0736_),
    .X(_0747_));
 sky130_fd_sc_hd__a211o_1 _1558_ (.A1(\MAC.add.b1[5] ),
    .A2(_0323_),
    .B1(_0728_),
    .C1(_0747_),
    .X(_0748_));
 sky130_fd_sc_hd__o31a_1 _1559_ (.A1(_0732_),
    .A2(_0742_),
    .A3(_0748_),
    .B1(\MAC.add.b1[15] ),
    .X(_0749_));
 sky130_fd_sc_hd__mux2_1 _1560_ (.A0(_0749_),
    .A1(\MAC.add.a1[15] ),
    .S(_0746_),
    .X(_0750_));
 sky130_fd_sc_hd__mux2_1 _1561_ (.A0(\MAC.add.b1[15] ),
    .A1(_0750_),
    .S(_0727_),
    .X(_0751_));
 sky130_fd_sc_hd__xnor2_1 _1562_ (.A(net29),
    .B(_0751_),
    .Y(_0752_));
 sky130_fd_sc_hd__nand2_1 _1563_ (.A(_0330_),
    .B(_0752_),
    .Y(_0753_));
 sky130_fd_sc_hd__a22o_1 _1564_ (.A1(_0665_),
    .A2(_0668_),
    .B1(_0753_),
    .B2(_0331_),
    .X(\MAC.add.c_add[15] ));
 sky130_fd_sc_hd__nand2_1 _1565_ (.A(\MAC.a[14] ),
    .B(\MAC.b[14] ),
    .Y(_0754_));
 sky130_fd_sc_hd__or2_1 _1566_ (.A(\MAC.a[14] ),
    .B(\MAC.b[14] ),
    .X(_0755_));
 sky130_fd_sc_hd__nand2_1 _1567_ (.A(_0754_),
    .B(_0755_),
    .Y(_0756_));
 sky130_fd_sc_hd__and2_1 _1568_ (.A(\MAC.a[12] ),
    .B(\MAC.b[12] ),
    .X(_0757_));
 sky130_fd_sc_hd__nor2_1 _1569_ (.A(\MAC.a[12] ),
    .B(\MAC.b[12] ),
    .Y(_0758_));
 sky130_fd_sc_hd__or2_1 _1570_ (.A(_0757_),
    .B(_0758_),
    .X(_0759_));
 sky130_fd_sc_hd__nand2_1 _1571_ (.A(\MAC.a[11] ),
    .B(\MAC.b[11] ),
    .Y(_0760_));
 sky130_fd_sc_hd__nand2_1 _1572_ (.A(\MAC.a[10] ),
    .B(\MAC.b[10] ),
    .Y(_0761_));
 sky130_fd_sc_hd__or2_1 _1573_ (.A(\MAC.a[10] ),
    .B(\MAC.b[10] ),
    .X(_0762_));
 sky130_fd_sc_hd__nand2_2 _1574_ (.A(_0761_),
    .B(_0762_),
    .Y(_0763_));
 sky130_fd_sc_hd__nand2_2 _1575_ (.A(\MAC.a[9] ),
    .B(\MAC.b[9] ),
    .Y(_0764_));
 sky130_fd_sc_hd__o21a_1 _1576_ (.A1(_0763_),
    .A2(_0764_),
    .B1(_0761_),
    .X(_0765_));
 sky130_fd_sc_hd__or2_1 _1577_ (.A(\MAC.a[11] ),
    .B(\MAC.b[11] ),
    .X(_0766_));
 sky130_fd_sc_hd__nand2_1 _1578_ (.A(_0760_),
    .B(_0766_),
    .Y(_0767_));
 sky130_fd_sc_hd__o21a_1 _1579_ (.A1(_0765_),
    .A2(_0767_),
    .B1(_0760_),
    .X(_0768_));
 sky130_fd_sc_hd__nor2_1 _1580_ (.A(_0759_),
    .B(_0768_),
    .Y(_0769_));
 sky130_fd_sc_hd__xor2_1 _1581_ (.A(\MAC.a[13] ),
    .B(\MAC.b[13] ),
    .X(_0770_));
 sky130_fd_sc_hd__xnor2_1 _1582_ (.A(\MAC.a[13] ),
    .B(\MAC.b[13] ),
    .Y(_0771_));
 sky130_fd_sc_hd__o21a_1 _1583_ (.A1(_0757_),
    .A2(_0769_),
    .B1(_0770_),
    .X(_0772_));
 sky130_fd_sc_hd__a21o_1 _1584_ (.A1(\MAC.a[13] ),
    .A2(\MAC.b[13] ),
    .B1(_0772_),
    .X(_0773_));
 sky130_fd_sc_hd__a21boi_1 _1585_ (.A1(_0755_),
    .A2(_0773_),
    .B1_N(_0754_),
    .Y(_0774_));
 sky130_fd_sc_hd__xor2_1 _1586_ (.A(_0756_),
    .B(_0773_),
    .X(_0775_));
 sky130_fd_sc_hd__or2_1 _1587_ (.A(\MAC.a[9] ),
    .B(\MAC.b[9] ),
    .X(_0776_));
 sky130_fd_sc_hd__nand2_2 _1588_ (.A(_0764_),
    .B(_0776_),
    .Y(_0777_));
 sky130_fd_sc_hd__nor2_1 _1589_ (.A(_0763_),
    .B(_0777_),
    .Y(_0778_));
 sky130_fd_sc_hd__or4_1 _1590_ (.A(_0759_),
    .B(_0763_),
    .C(_0767_),
    .D(_0777_),
    .X(_0779_));
 sky130_fd_sc_hd__or2_1 _1591_ (.A(_0771_),
    .B(_0779_),
    .X(_0780_));
 sky130_fd_sc_hd__xnor2_1 _1592_ (.A(_0775_),
    .B(_0780_),
    .Y(_0781_));
 sky130_fd_sc_hd__or2_1 _1593_ (.A(_0774_),
    .B(_0781_),
    .X(_0782_));
 sky130_fd_sc_hd__or2_1 _1594_ (.A(_0755_),
    .B(_0773_),
    .X(_0783_));
 sky130_fd_sc_hd__nand2_1 _1595_ (.A(_0782_),
    .B(net25),
    .Y(_0784_));
 sky130_fd_sc_hd__nor3_1 _1596_ (.A(_0757_),
    .B(_0769_),
    .C(_0770_),
    .Y(_0785_));
 sky130_fd_sc_hd__nor2_1 _1597_ (.A(_0772_),
    .B(_0785_),
    .Y(_0786_));
 sky130_fd_sc_hd__and2_1 _1598_ (.A(_0759_),
    .B(_0768_),
    .X(_0787_));
 sky130_fd_sc_hd__nor2_1 _1599_ (.A(_0769_),
    .B(_0787_),
    .Y(_0788_));
 sky130_fd_sc_hd__xor2_1 _1600_ (.A(_0765_),
    .B(_0767_),
    .X(_0789_));
 sky130_fd_sc_hd__nand2_1 _1601_ (.A(_0778_),
    .B(_0789_),
    .Y(_0790_));
 sky130_fd_sc_hd__or2_1 _1602_ (.A(_0778_),
    .B(_0789_),
    .X(_0791_));
 sky130_fd_sc_hd__and2_1 _1603_ (.A(_0790_),
    .B(_0791_),
    .X(_0792_));
 sky130_fd_sc_hd__xor2_2 _1604_ (.A(_0763_),
    .B(_0764_),
    .X(_0793_));
 sky130_fd_sc_hd__and3_1 _1605_ (.A(_0777_),
    .B(_0789_),
    .C(_0793_),
    .X(_0794_));
 sky130_fd_sc_hd__and4b_1 _1606_ (.A_N(_0774_),
    .B(_0786_),
    .C(_0788_),
    .D(_0794_),
    .X(_0795_));
 sky130_fd_sc_hd__nand2_2 _1607_ (.A(net59),
    .B(net57),
    .Y(_0796_));
 sky130_fd_sc_hd__nand2_1 _1608_ (.A(net44),
    .B(net41),
    .Y(_0797_));
 sky130_fd_sc_hd__and2_1 _1609_ (.A(net68),
    .B(net66),
    .X(_0798_));
 sky130_fd_sc_hd__nand2_1 _1610_ (.A(net68),
    .B(net66),
    .Y(_0799_));
 sky130_fd_sc_hd__and2_1 _1611_ (.A(net75),
    .B(net74),
    .X(_0800_));
 sky130_fd_sc_hd__nand2_1 _1612_ (.A(net63),
    .B(net61),
    .Y(_0801_));
 sky130_fd_sc_hd__and4_1 _1613_ (.A(net46),
    .B(\MAC.a[7] ),
    .C(net42),
    .D(\MAC.a[15] ),
    .X(_0802_));
 sky130_fd_sc_hd__and4_1 _1614_ (.A(\MAC.a[14] ),
    .B(\MAC.a[13] ),
    .C(net50),
    .D(net48),
    .X(_0803_));
 sky130_fd_sc_hd__and4_1 _1615_ (.A(\MAC.a[10] ),
    .B(\MAC.a[9] ),
    .C(\MAC.a[12] ),
    .D(\MAC.a[11] ),
    .X(_0804_));
 sky130_fd_sc_hd__and4_1 _1616_ (.A(net59),
    .B(net57),
    .C(net54),
    .D(net52),
    .X(_0805_));
 sky130_fd_sc_hd__and4_1 _1617_ (.A(\MAC.b[10] ),
    .B(\MAC.b[9] ),
    .C(\MAC.b[12] ),
    .D(\MAC.b[11] ),
    .X(_0806_));
 sky130_fd_sc_hd__and3_1 _1618_ (.A(_0798_),
    .B(_0800_),
    .C(_0806_),
    .X(_0807_));
 sky130_fd_sc_hd__and4_1 _1619_ (.A(net65),
    .B(net63),
    .C(net61),
    .D(\MAC.b[15] ),
    .X(_0808_));
 sky130_fd_sc_hd__and4_1 _1620_ (.A(_0802_),
    .B(_0803_),
    .C(_0804_),
    .D(_0805_),
    .X(_0809_));
 sky130_fd_sc_hd__and4_1 _1621_ (.A(\MAC.b[14] ),
    .B(\MAC.b[13] ),
    .C(\MAC.b[2] ),
    .D(\MAC.b[3] ),
    .X(_0810_));
 sky130_fd_sc_hd__a31o_1 _1622_ (.A1(_0807_),
    .A2(_0808_),
    .A3(_0810_),
    .B1(_0809_),
    .X(_0811_));
 sky130_fd_sc_hd__a21oi_1 _1623_ (.A1(_0775_),
    .A2(_0795_),
    .B1(_0811_),
    .Y(_0812_));
 sky130_fd_sc_hd__and2_1 _1624_ (.A(net41),
    .B(net60),
    .X(_0813_));
 sky130_fd_sc_hd__nor2_1 _1625_ (.A(net41),
    .B(net60),
    .Y(_0814_));
 sky130_fd_sc_hd__or2_1 _1626_ (.A(_0813_),
    .B(_0814_),
    .X(_0815_));
 sky130_fd_sc_hd__nand2_1 _1627_ (.A(net44),
    .B(net62),
    .Y(_0816_));
 sky130_fd_sc_hd__o21bai_2 _1628_ (.A1(_0814_),
    .A2(_0816_),
    .B1_N(_0813_),
    .Y(_0817_));
 sky130_fd_sc_hd__nand2_1 _1629_ (.A(net46),
    .B(net61),
    .Y(_0818_));
 sky130_fd_sc_hd__nor2_1 _1630_ (.A(_0816_),
    .B(_0818_),
    .Y(_0819_));
 sky130_fd_sc_hd__nand2_1 _1631_ (.A(_0816_),
    .B(_0818_),
    .Y(_0820_));
 sky130_fd_sc_hd__and2b_1 _1632_ (.A_N(_0819_),
    .B(_0820_),
    .X(_0821_));
 sky130_fd_sc_hd__nand2_1 _1633_ (.A(net41),
    .B(net65),
    .Y(_0822_));
 sky130_fd_sc_hd__a31o_1 _1634_ (.A1(net41),
    .A2(net65),
    .A3(_0820_),
    .B1(_0819_),
    .X(_0823_));
 sky130_fd_sc_hd__or2_1 _1635_ (.A(_0797_),
    .B(_0801_),
    .X(_0824_));
 sky130_fd_sc_hd__a22o_1 _1636_ (.A1(net41),
    .A2(net63),
    .B1(net60),
    .B2(net44),
    .X(_0825_));
 sky130_fd_sc_hd__and3_1 _1637_ (.A(net65),
    .B(_0824_),
    .C(_0825_),
    .X(_0826_));
 sky130_fd_sc_hd__a21oi_1 _1638_ (.A1(_0824_),
    .A2(_0825_),
    .B1(net65),
    .Y(_0827_));
 sky130_fd_sc_hd__nor2_1 _1639_ (.A(_0826_),
    .B(_0827_),
    .Y(_0828_));
 sky130_fd_sc_hd__and2_1 _1640_ (.A(net46),
    .B(_0828_),
    .X(_0829_));
 sky130_fd_sc_hd__inv_2 _1641_ (.A(_0829_),
    .Y(_0830_));
 sky130_fd_sc_hd__xnor2_1 _1642_ (.A(net46),
    .B(_0828_),
    .Y(_0831_));
 sky130_fd_sc_hd__xnor2_1 _1643_ (.A(_0821_),
    .B(_0822_),
    .Y(_0832_));
 sky130_fd_sc_hd__nand2_1 _1644_ (.A(net48),
    .B(_0832_),
    .Y(_0833_));
 sky130_fd_sc_hd__nor2_1 _1645_ (.A(_0831_),
    .B(_0833_),
    .Y(_0834_));
 sky130_fd_sc_hd__and2_1 _1646_ (.A(_0831_),
    .B(_0833_),
    .X(_0835_));
 sky130_fd_sc_hd__nor2_1 _1647_ (.A(_0834_),
    .B(_0835_),
    .Y(_0836_));
 sky130_fd_sc_hd__and2_1 _1648_ (.A(_0823_),
    .B(_0836_),
    .X(_0837_));
 sky130_fd_sc_hd__nor2_1 _1649_ (.A(_0823_),
    .B(_0836_),
    .Y(_0838_));
 sky130_fd_sc_hd__or2_1 _1650_ (.A(_0837_),
    .B(_0838_),
    .X(_0839_));
 sky130_fd_sc_hd__or2_1 _1651_ (.A(net48),
    .B(_0832_),
    .X(_0840_));
 sky130_fd_sc_hd__nand2_1 _1652_ (.A(_0833_),
    .B(_0840_),
    .Y(_0841_));
 sky130_fd_sc_hd__a22o_1 _1653_ (.A1(\MAC.a[6] ),
    .A2(net62),
    .B1(net60),
    .B2(net48),
    .X(_0842_));
 sky130_fd_sc_hd__nand2_1 _1654_ (.A(net48),
    .B(net62),
    .Y(_0843_));
 sky130_fd_sc_hd__nor2_1 _1655_ (.A(_0818_),
    .B(_0843_),
    .Y(_0844_));
 sky130_fd_sc_hd__o21a_1 _1656_ (.A1(_0818_),
    .A2(_0843_),
    .B1(_0842_),
    .X(_0845_));
 sky130_fd_sc_hd__nand2_1 _1657_ (.A(\MAC.a[7] ),
    .B(net65),
    .Y(_0846_));
 sky130_fd_sc_hd__xnor2_1 _1658_ (.A(_0845_),
    .B(_0846_),
    .Y(_0847_));
 sky130_fd_sc_hd__nand2_1 _1659_ (.A(net49),
    .B(_0847_),
    .Y(_0848_));
 sky130_fd_sc_hd__xor2_1 _1660_ (.A(_0841_),
    .B(_0848_),
    .X(_0849_));
 sky130_fd_sc_hd__a31oi_1 _1661_ (.A1(\MAC.a[7] ),
    .A2(net65),
    .A3(_0842_),
    .B1(_0844_),
    .Y(_0850_));
 sky130_fd_sc_hd__nand2_1 _1662_ (.A(net41),
    .B(net68),
    .Y(_0851_));
 sky130_fd_sc_hd__a21o_1 _1663_ (.A1(net66),
    .A2(_0851_),
    .B1(_0850_),
    .X(_0852_));
 sky130_fd_sc_hd__nand2_1 _1664_ (.A(_0850_),
    .B(_0851_),
    .Y(_0853_));
 sky130_fd_sc_hd__o21ai_1 _1665_ (.A1(_0329_),
    .A2(_0853_),
    .B1(_0852_),
    .Y(_0854_));
 sky130_fd_sc_hd__nand2_1 _1666_ (.A(_0849_),
    .B(_0854_),
    .Y(_0855_));
 sky130_fd_sc_hd__o21a_1 _1667_ (.A1(_0841_),
    .A2(_0848_),
    .B1(_0855_),
    .X(_0856_));
 sky130_fd_sc_hd__nor2_1 _1668_ (.A(_0839_),
    .B(_0856_),
    .Y(_0857_));
 sky130_fd_sc_hd__and2_1 _1669_ (.A(_0839_),
    .B(_0856_),
    .X(_0858_));
 sky130_fd_sc_hd__nor2_1 _1670_ (.A(_0857_),
    .B(_0858_),
    .Y(_0859_));
 sky130_fd_sc_hd__and3_1 _1671_ (.A(net66),
    .B(_0853_),
    .C(_0859_),
    .X(_0860_));
 sky130_fd_sc_hd__a21oi_1 _1672_ (.A1(net66),
    .A2(_0853_),
    .B1(_0859_),
    .Y(_0861_));
 sky130_fd_sc_hd__or2_1 _1673_ (.A(_0860_),
    .B(_0861_),
    .X(_0862_));
 sky130_fd_sc_hd__or2_1 _1674_ (.A(_0849_),
    .B(_0854_),
    .X(_0863_));
 sky130_fd_sc_hd__and2_1 _1675_ (.A(_0855_),
    .B(_0863_),
    .X(_0864_));
 sky130_fd_sc_hd__or2_1 _1676_ (.A(net49),
    .B(_0847_),
    .X(_0865_));
 sky130_fd_sc_hd__nand2_1 _1677_ (.A(_0848_),
    .B(_0865_),
    .Y(_0866_));
 sky130_fd_sc_hd__nand2_1 _1678_ (.A(net49),
    .B(net60),
    .Y(_0867_));
 sky130_fd_sc_hd__nor2_1 _1679_ (.A(_0843_),
    .B(_0867_),
    .Y(_0868_));
 sky130_fd_sc_hd__xor2_1 _1680_ (.A(_0843_),
    .B(_0867_),
    .X(_0869_));
 sky130_fd_sc_hd__nand2_1 _1681_ (.A(net45),
    .B(net64),
    .Y(_0870_));
 sky130_fd_sc_hd__xnor2_1 _1682_ (.A(_0869_),
    .B(_0870_),
    .Y(_0871_));
 sky130_fd_sc_hd__nand2_1 _1683_ (.A(net53),
    .B(_0871_),
    .Y(_0872_));
 sky130_fd_sc_hd__a31o_1 _1684_ (.A1(net46),
    .A2(net64),
    .A3(_0869_),
    .B1(_0868_),
    .X(_0873_));
 sky130_fd_sc_hd__or2_1 _1685_ (.A(\MAC.b[4] ),
    .B(\MAC.b[5] ),
    .X(_0874_));
 sky130_fd_sc_hd__and2b_1 _1686_ (.A_N(net41),
    .B(net68),
    .X(_0875_));
 sky130_fd_sc_hd__a31o_1 _1687_ (.A1(net41),
    .A2(_0799_),
    .A3(_0874_),
    .B1(_0875_),
    .X(_0876_));
 sky130_fd_sc_hd__xor2_1 _1688_ (.A(_0873_),
    .B(_0876_),
    .X(_0877_));
 sky130_fd_sc_hd__a22o_1 _1689_ (.A1(net41),
    .A2(net68),
    .B1(net66),
    .B2(net44),
    .X(_0878_));
 sky130_fd_sc_hd__o21a_1 _1690_ (.A1(_0797_),
    .A2(_0799_),
    .B1(_0878_),
    .X(_0879_));
 sky130_fd_sc_hd__o2bb2a_1 _1691_ (.A1_N(net71),
    .A2_N(_0878_),
    .B1(_0799_),
    .B2(_0797_),
    .X(_0880_));
 sky130_fd_sc_hd__nand2b_1 _1692_ (.A_N(_0880_),
    .B(_0877_),
    .Y(_0881_));
 sky130_fd_sc_hd__xnor2_1 _1693_ (.A(_0877_),
    .B(_0880_),
    .Y(_0882_));
 sky130_fd_sc_hd__xor2_1 _1694_ (.A(_0866_),
    .B(_0872_),
    .X(_0883_));
 sky130_fd_sc_hd__and2_1 _1695_ (.A(_0882_),
    .B(_0883_),
    .X(_0884_));
 sky130_fd_sc_hd__o21ba_1 _1696_ (.A1(_0866_),
    .A2(_0872_),
    .B1_N(_0884_),
    .X(_0885_));
 sky130_fd_sc_hd__nand2b_1 _1697_ (.A_N(_0885_),
    .B(_0864_),
    .Y(_0886_));
 sky130_fd_sc_hd__a21bo_1 _1698_ (.A1(_0873_),
    .A2(_0876_),
    .B1_N(_0881_),
    .X(_0887_));
 sky130_fd_sc_hd__xnor2_1 _1699_ (.A(_0864_),
    .B(_0885_),
    .Y(_0888_));
 sky130_fd_sc_hd__nand2_1 _1700_ (.A(_0887_),
    .B(_0888_),
    .Y(_0889_));
 sky130_fd_sc_hd__a21oi_1 _1701_ (.A1(_0886_),
    .A2(_0889_),
    .B1(_0862_),
    .Y(_0890_));
 sky130_fd_sc_hd__o21ba_1 _1702_ (.A1(_0797_),
    .A2(_0801_),
    .B1_N(_0826_),
    .X(_0891_));
 sky130_fd_sc_hd__nand2_1 _1703_ (.A(net63),
    .B(_0813_),
    .Y(_0892_));
 sky130_fd_sc_hd__or2_1 _1704_ (.A(net63),
    .B(_0813_),
    .X(_0893_));
 sky130_fd_sc_hd__and3_1 _1705_ (.A(net44),
    .B(_0892_),
    .C(_0893_),
    .X(_0894_));
 sky130_fd_sc_hd__a21oi_1 _1706_ (.A1(_0892_),
    .A2(_0893_),
    .B1(net44),
    .Y(_0895_));
 sky130_fd_sc_hd__or2_1 _1707_ (.A(_0894_),
    .B(_0895_),
    .X(_0896_));
 sky130_fd_sc_hd__nor2_1 _1708_ (.A(_0830_),
    .B(_0896_),
    .Y(_0897_));
 sky130_fd_sc_hd__and2_1 _1709_ (.A(_0830_),
    .B(_0896_),
    .X(_0898_));
 sky130_fd_sc_hd__nor2_1 _1710_ (.A(_0897_),
    .B(_0898_),
    .Y(_0899_));
 sky130_fd_sc_hd__and2b_1 _1711_ (.A_N(_0891_),
    .B(_0899_),
    .X(_0900_));
 sky130_fd_sc_hd__xnor2_1 _1712_ (.A(_0891_),
    .B(_0899_),
    .Y(_0901_));
 sky130_fd_sc_hd__o21ai_1 _1713_ (.A1(_0834_),
    .A2(_0837_),
    .B1(_0901_),
    .Y(_0902_));
 sky130_fd_sc_hd__or3_1 _1714_ (.A(_0834_),
    .B(_0837_),
    .C(_0901_),
    .X(_0903_));
 sky130_fd_sc_hd__and2_1 _1715_ (.A(_0902_),
    .B(_0903_),
    .X(_0904_));
 sky130_fd_sc_hd__o21ai_1 _1716_ (.A1(_0857_),
    .A2(_0860_),
    .B1(_0904_),
    .Y(_0905_));
 sky130_fd_sc_hd__or3_1 _1717_ (.A(_0857_),
    .B(_0860_),
    .C(_0904_),
    .X(_0906_));
 sky130_fd_sc_hd__and2_1 _1718_ (.A(_0905_),
    .B(_0906_),
    .X(_0907_));
 sky130_fd_sc_hd__nand2_1 _1719_ (.A(_0890_),
    .B(_0907_),
    .Y(_0908_));
 sky130_fd_sc_hd__and3_1 _1720_ (.A(_0862_),
    .B(_0886_),
    .C(_0889_),
    .X(_0909_));
 sky130_fd_sc_hd__or2_1 _1721_ (.A(_0887_),
    .B(_0888_),
    .X(_0910_));
 sky130_fd_sc_hd__nand2_1 _1722_ (.A(_0889_),
    .B(_0910_),
    .Y(_0911_));
 sky130_fd_sc_hd__nor2_1 _1723_ (.A(_0882_),
    .B(_0883_),
    .Y(_0912_));
 sky130_fd_sc_hd__or2_1 _1724_ (.A(_0884_),
    .B(_0912_),
    .X(_0913_));
 sky130_fd_sc_hd__or2_1 _1725_ (.A(net53),
    .B(_0871_),
    .X(_0914_));
 sky130_fd_sc_hd__nand2_1 _1726_ (.A(_0872_),
    .B(_0914_),
    .Y(_0915_));
 sky130_fd_sc_hd__and3_1 _1727_ (.A(net57),
    .B(\MAC.a[2] ),
    .C(net74),
    .X(_0916_));
 sky130_fd_sc_hd__nand3_1 _1728_ (.A(net56),
    .B(net55),
    .C(net73),
    .Y(_0917_));
 sky130_fd_sc_hd__nand2_1 _1729_ (.A(net51),
    .B(net62),
    .Y(_0918_));
 sky130_fd_sc_hd__or2_1 _1730_ (.A(_0867_),
    .B(_0918_),
    .X(_0919_));
 sky130_fd_sc_hd__a22o_1 _1731_ (.A1(net49),
    .A2(net62),
    .B1(net60),
    .B2(net51),
    .X(_0920_));
 sky130_fd_sc_hd__nand2_1 _1732_ (.A(_0919_),
    .B(_0920_),
    .Y(_0921_));
 sky130_fd_sc_hd__nand2_1 _1733_ (.A(net47),
    .B(net64),
    .Y(_0922_));
 sky130_fd_sc_hd__xnor2_1 _1734_ (.A(_0921_),
    .B(_0922_),
    .Y(_0923_));
 sky130_fd_sc_hd__a21o_1 _1735_ (.A1(net56),
    .A2(net73),
    .B1(net55),
    .X(_0924_));
 sky130_fd_sc_hd__nand2_1 _1736_ (.A(_0917_),
    .B(_0924_),
    .Y(_0925_));
 sky130_fd_sc_hd__or2_1 _1737_ (.A(_0923_),
    .B(_0925_),
    .X(_0926_));
 sky130_fd_sc_hd__a21o_1 _1738_ (.A1(_0917_),
    .A2(_0926_),
    .B1(_0915_),
    .X(_0927_));
 sky130_fd_sc_hd__o21ai_1 _1739_ (.A1(_0921_),
    .A2(_0922_),
    .B1(_0919_),
    .Y(_0928_));
 sky130_fd_sc_hd__xnor2_1 _1740_ (.A(net70),
    .B(_0879_),
    .Y(_0929_));
 sky130_fd_sc_hd__nand2b_1 _1741_ (.A_N(_0929_),
    .B(_0928_),
    .Y(_0930_));
 sky130_fd_sc_hd__xnor2_1 _1742_ (.A(_0928_),
    .B(_0929_),
    .Y(_0931_));
 sky130_fd_sc_hd__and4_1 _1743_ (.A(net45),
    .B(net43),
    .C(net69),
    .D(net67),
    .X(_0932_));
 sky130_fd_sc_hd__a22oi_1 _1744_ (.A1(net43),
    .A2(net69),
    .B1(net67),
    .B2(net45),
    .Y(_0933_));
 sky130_fd_sc_hd__and4bb_1 _1745_ (.A_N(_0932_),
    .B_N(_0933_),
    .C(net42),
    .D(net70),
    .X(_0934_));
 sky130_fd_sc_hd__or2_1 _1746_ (.A(_0932_),
    .B(_0934_),
    .X(_0935_));
 sky130_fd_sc_hd__xnor2_1 _1747_ (.A(_0931_),
    .B(_0935_),
    .Y(_0936_));
 sky130_fd_sc_hd__nand3_1 _1748_ (.A(_0915_),
    .B(_0917_),
    .C(_0926_),
    .Y(_0937_));
 sky130_fd_sc_hd__nand2_1 _1749_ (.A(_0927_),
    .B(_0937_),
    .Y(_0938_));
 sky130_fd_sc_hd__or2_1 _1750_ (.A(_0936_),
    .B(_0938_),
    .X(_0939_));
 sky130_fd_sc_hd__a21oi_1 _1751_ (.A1(_0927_),
    .A2(_0939_),
    .B1(_0913_),
    .Y(_0940_));
 sky130_fd_sc_hd__a21bo_1 _1752_ (.A1(_0931_),
    .A2(_0935_),
    .B1_N(_0930_),
    .X(_0941_));
 sky130_fd_sc_hd__and3_1 _1753_ (.A(_0913_),
    .B(_0927_),
    .C(_0939_),
    .X(_0942_));
 sky130_fd_sc_hd__nor2_1 _1754_ (.A(_0940_),
    .B(_0942_),
    .Y(_0943_));
 sky130_fd_sc_hd__a21oi_1 _1755_ (.A1(_0941_),
    .A2(_0943_),
    .B1(_0940_),
    .Y(_0944_));
 sky130_fd_sc_hd__or2_1 _1756_ (.A(_0911_),
    .B(_0944_),
    .X(_0945_));
 sky130_fd_sc_hd__or3_1 _1757_ (.A(_0890_),
    .B(_0909_),
    .C(_0945_),
    .X(_0946_));
 sky130_fd_sc_hd__o21ai_1 _1758_ (.A1(_0890_),
    .A2(_0909_),
    .B1(_0945_),
    .Y(_0947_));
 sky130_fd_sc_hd__and2_1 _1759_ (.A(_0946_),
    .B(_0947_),
    .X(_0948_));
 sky130_fd_sc_hd__xnor2_1 _1760_ (.A(_0911_),
    .B(_0944_),
    .Y(_0949_));
 sky130_fd_sc_hd__xor2_1 _1761_ (.A(_0941_),
    .B(_0943_),
    .X(_0950_));
 sky130_fd_sc_hd__nand2_1 _1762_ (.A(_0936_),
    .B(_0938_),
    .Y(_0951_));
 sky130_fd_sc_hd__xnor2_1 _1763_ (.A(_0923_),
    .B(_0925_),
    .Y(_0952_));
 sky130_fd_sc_hd__xnor2_1 _1764_ (.A(net56),
    .B(net73),
    .Y(_0953_));
 sky130_fd_sc_hd__and3_1 _1765_ (.A(net42),
    .B(net76),
    .C(net73),
    .X(_0954_));
 sky130_fd_sc_hd__a21o_1 _1766_ (.A1(net42),
    .A2(net73),
    .B1(net76),
    .X(_0955_));
 sky130_fd_sc_hd__o21ai_1 _1767_ (.A1(net58),
    .A2(_0954_),
    .B1(_0955_),
    .Y(_0956_));
 sky130_fd_sc_hd__xor2_1 _1768_ (.A(_0953_),
    .B(_0956_),
    .X(_0957_));
 sky130_fd_sc_hd__and4_1 _1769_ (.A(net55),
    .B(net51),
    .C(net62),
    .D(net60),
    .X(_0958_));
 sky130_fd_sc_hd__nand2_1 _1770_ (.A(net55),
    .B(net60),
    .Y(_0959_));
 sky130_fd_sc_hd__a21o_1 _1771_ (.A1(_0918_),
    .A2(_0959_),
    .B1(_0958_),
    .X(_0960_));
 sky130_fd_sc_hd__nand2_1 _1772_ (.A(net49),
    .B(net64),
    .Y(_0961_));
 sky130_fd_sc_hd__xor2_1 _1773_ (.A(_0960_),
    .B(_0961_),
    .X(_0962_));
 sky130_fd_sc_hd__nand2_1 _1774_ (.A(_0957_),
    .B(_0962_),
    .Y(_0963_));
 sky130_fd_sc_hd__o21ai_1 _1775_ (.A1(_0953_),
    .A2(_0956_),
    .B1(_0963_),
    .Y(_0964_));
 sky130_fd_sc_hd__and2b_1 _1776_ (.A_N(_0952_),
    .B(_0964_),
    .X(_0965_));
 sky130_fd_sc_hd__o21ba_1 _1777_ (.A1(_0960_),
    .A2(_0961_),
    .B1_N(_0958_),
    .X(_0966_));
 sky130_fd_sc_hd__o2bb2a_1 _1778_ (.A1_N(net42),
    .A2_N(net70),
    .B1(_0932_),
    .B2(_0933_),
    .X(_0967_));
 sky130_fd_sc_hd__nor2_1 _1779_ (.A(_0934_),
    .B(_0967_),
    .Y(_0968_));
 sky130_fd_sc_hd__or3_1 _1780_ (.A(_0934_),
    .B(_0966_),
    .C(_0967_),
    .X(_0969_));
 sky130_fd_sc_hd__xnor2_1 _1781_ (.A(_0966_),
    .B(_0968_),
    .Y(_0970_));
 sky130_fd_sc_hd__and4_1 _1782_ (.A(net47),
    .B(net45),
    .C(net69),
    .D(net67),
    .X(_0971_));
 sky130_fd_sc_hd__a22o_1 _1783_ (.A1(net45),
    .A2(net69),
    .B1(net67),
    .B2(net47),
    .X(_0972_));
 sky130_fd_sc_hd__and2b_1 _1784_ (.A_N(_0971_),
    .B(_0972_),
    .X(_0973_));
 sky130_fd_sc_hd__nand2_1 _1785_ (.A(net43),
    .B(net70),
    .Y(_0974_));
 sky130_fd_sc_hd__a31oi_1 _1786_ (.A1(net43),
    .A2(net70),
    .A3(_0972_),
    .B1(_0971_),
    .Y(_0975_));
 sky130_fd_sc_hd__nand2b_1 _1787_ (.A_N(_0975_),
    .B(_0970_),
    .Y(_0976_));
 sky130_fd_sc_hd__xor2_1 _1788_ (.A(_0970_),
    .B(_0975_),
    .X(_0977_));
 sky130_fd_sc_hd__xor2_1 _1789_ (.A(_0952_),
    .B(_0964_),
    .X(_0978_));
 sky130_fd_sc_hd__nor2_1 _1790_ (.A(_0977_),
    .B(_0978_),
    .Y(_0979_));
 sky130_fd_sc_hd__o211a_1 _1791_ (.A1(_0965_),
    .A2(_0979_),
    .B1(_0939_),
    .C1(_0951_),
    .X(_0980_));
 sky130_fd_sc_hd__a211oi_1 _1792_ (.A1(_0939_),
    .A2(_0951_),
    .B1(_0965_),
    .C1(_0979_),
    .Y(_0981_));
 sky130_fd_sc_hd__a211oi_1 _1793_ (.A1(_0969_),
    .A2(_0976_),
    .B1(_0980_),
    .C1(_0981_),
    .Y(_0982_));
 sky130_fd_sc_hd__o21a_1 _1794_ (.A1(_0980_),
    .A2(_0982_),
    .B1(_0950_),
    .X(_0983_));
 sky130_fd_sc_hd__and2b_1 _1795_ (.A_N(_0949_),
    .B(_0983_),
    .X(_0984_));
 sky130_fd_sc_hd__xnor2_1 _1796_ (.A(_0949_),
    .B(_0983_),
    .Y(_0985_));
 sky130_fd_sc_hd__or3_1 _1797_ (.A(_0950_),
    .B(_0980_),
    .C(_0982_),
    .X(_0986_));
 sky130_fd_sc_hd__and2b_1 _1798_ (.A_N(_0983_),
    .B(_0986_),
    .X(_0987_));
 sky130_fd_sc_hd__o211a_1 _1799_ (.A1(_0980_),
    .A2(_0981_),
    .B1(_0969_),
    .C1(_0976_),
    .X(_0988_));
 sky130_fd_sc_hd__nor2_1 _1800_ (.A(_0982_),
    .B(_0988_),
    .Y(_0989_));
 sky130_fd_sc_hd__and2_1 _1801_ (.A(_0977_),
    .B(_0978_),
    .X(_0990_));
 sky130_fd_sc_hd__or2_1 _1802_ (.A(_0957_),
    .B(_0962_),
    .X(_0991_));
 sky130_fd_sc_hd__nand2_1 _1803_ (.A(_0963_),
    .B(_0991_),
    .Y(_0992_));
 sky130_fd_sc_hd__and4_1 _1804_ (.A(net56),
    .B(net55),
    .C(net62),
    .D(net60),
    .X(_0993_));
 sky130_fd_sc_hd__a22o_1 _1805_ (.A1(net55),
    .A2(net62),
    .B1(net60),
    .B2(net56),
    .X(_0994_));
 sky130_fd_sc_hd__nand2b_1 _1806_ (.A_N(_0993_),
    .B(_0994_),
    .Y(_0995_));
 sky130_fd_sc_hd__nand2_1 _1807_ (.A(net51),
    .B(net64),
    .Y(_0996_));
 sky130_fd_sc_hd__xnor2_1 _1808_ (.A(_0995_),
    .B(_0996_),
    .Y(_0997_));
 sky130_fd_sc_hd__a21boi_1 _1809_ (.A1(_0328_),
    .A2(_0954_),
    .B1_N(_0955_),
    .Y(_0998_));
 sky130_fd_sc_hd__xnor2_1 _1810_ (.A(net58),
    .B(_0998_),
    .Y(_0999_));
 sky130_fd_sc_hd__nor2_1 _1811_ (.A(_0997_),
    .B(_0999_),
    .Y(_1000_));
 sky130_fd_sc_hd__a41o_1 _1812_ (.A1(net58),
    .A2(net43),
    .A3(net42),
    .A4(_0800_),
    .B1(_1000_),
    .X(_1001_));
 sky130_fd_sc_hd__nand2b_1 _1813_ (.A_N(_0992_),
    .B(_1001_),
    .Y(_1002_));
 sky130_fd_sc_hd__xnor2_1 _1814_ (.A(_0992_),
    .B(_1001_),
    .Y(_1003_));
 sky130_fd_sc_hd__and4_1 _1815_ (.A(net49),
    .B(net47),
    .C(net69),
    .D(net67),
    .X(_1004_));
 sky130_fd_sc_hd__a22o_1 _1816_ (.A1(net47),
    .A2(net69),
    .B1(net67),
    .B2(net49),
    .X(_1005_));
 sky130_fd_sc_hd__and2b_1 _1817_ (.A_N(_1004_),
    .B(_1005_),
    .X(_1006_));
 sky130_fd_sc_hd__nand2_1 _1818_ (.A(net45),
    .B(net70),
    .Y(_1007_));
 sky130_fd_sc_hd__a31oi_2 _1819_ (.A1(net45),
    .A2(net70),
    .A3(_1005_),
    .B1(_1004_),
    .Y(_1008_));
 sky130_fd_sc_hd__a31o_1 _1820_ (.A1(net51),
    .A2(net64),
    .A3(_0994_),
    .B1(_0993_),
    .X(_1009_));
 sky130_fd_sc_hd__xnor2_1 _1821_ (.A(_0973_),
    .B(_0974_),
    .Y(_1010_));
 sky130_fd_sc_hd__and2_1 _1822_ (.A(_1009_),
    .B(_1010_),
    .X(_1011_));
 sky130_fd_sc_hd__nor2_1 _1823_ (.A(_1009_),
    .B(_1010_),
    .Y(_1012_));
 sky130_fd_sc_hd__nor2_1 _1824_ (.A(_1011_),
    .B(_1012_),
    .Y(_1013_));
 sky130_fd_sc_hd__and2b_1 _1825_ (.A_N(_1008_),
    .B(_1013_),
    .X(_1014_));
 sky130_fd_sc_hd__xnor2_1 _1826_ (.A(_1008_),
    .B(_1013_),
    .Y(_1015_));
 sky130_fd_sc_hd__nand2_1 _1827_ (.A(_1003_),
    .B(_1015_),
    .Y(_1016_));
 sky130_fd_sc_hd__a211o_1 _1828_ (.A1(_1002_),
    .A2(_1016_),
    .B1(_0979_),
    .C1(_0990_),
    .X(_1017_));
 sky130_fd_sc_hd__inv_2 _1829_ (.A(_1017_),
    .Y(_1018_));
 sky130_fd_sc_hd__o211ai_1 _1830_ (.A1(_0979_),
    .A2(_0990_),
    .B1(_1002_),
    .C1(_1016_),
    .Y(_1019_));
 sky130_fd_sc_hd__o211a_1 _1831_ (.A1(_1011_),
    .A2(_1014_),
    .B1(_1017_),
    .C1(_1019_),
    .X(_1020_));
 sky130_fd_sc_hd__nor2_1 _1832_ (.A(_1018_),
    .B(_1020_),
    .Y(_1021_));
 sky130_fd_sc_hd__and2b_1 _1833_ (.A_N(_1021_),
    .B(_0989_),
    .X(_1022_));
 sky130_fd_sc_hd__and2_1 _1834_ (.A(_0987_),
    .B(_1022_),
    .X(_1023_));
 sky130_fd_sc_hd__nor2_1 _1835_ (.A(_0987_),
    .B(_1022_),
    .Y(_1024_));
 sky130_fd_sc_hd__or2_1 _1836_ (.A(_1023_),
    .B(_1024_),
    .X(_1025_));
 sky130_fd_sc_hd__xnor2_1 _1837_ (.A(_0989_),
    .B(_1021_),
    .Y(_1026_));
 sky130_fd_sc_hd__a211oi_1 _1838_ (.A1(_1017_),
    .A2(_1019_),
    .B1(_1011_),
    .C1(_1014_),
    .Y(_1027_));
 sky130_fd_sc_hd__xnor2_1 _1839_ (.A(_1003_),
    .B(_1015_),
    .Y(_1028_));
 sky130_fd_sc_hd__and2_1 _1840_ (.A(_0997_),
    .B(_0999_),
    .X(_1029_));
 sky130_fd_sc_hd__or2_1 _1841_ (.A(_1000_),
    .B(_1029_),
    .X(_1030_));
 sky130_fd_sc_hd__a22oi_1 _1842_ (.A1(net42),
    .A2(net76),
    .B1(net73),
    .B2(net44),
    .Y(_1031_));
 sky130_fd_sc_hd__a31o_1 _1843_ (.A1(net43),
    .A2(net42),
    .A3(_0800_),
    .B1(_1031_),
    .X(_1032_));
 sky130_fd_sc_hd__nand2_1 _1844_ (.A(net46),
    .B(net75),
    .Y(_1033_));
 sky130_fd_sc_hd__nand2_1 _1845_ (.A(net43),
    .B(net76),
    .Y(_1034_));
 sky130_fd_sc_hd__and4_1 _1846_ (.A(net45),
    .B(net44),
    .C(net76),
    .D(net73),
    .X(_1035_));
 sky130_fd_sc_hd__nand2b_1 _1847_ (.A_N(_1032_),
    .B(_1035_),
    .Y(_1036_));
 sky130_fd_sc_hd__nor2_1 _1848_ (.A(_0796_),
    .B(_0801_),
    .Y(_1037_));
 sky130_fd_sc_hd__a22o_1 _1849_ (.A1(net57),
    .A2(net63),
    .B1(net61),
    .B2(net58),
    .X(_1038_));
 sky130_fd_sc_hd__o21a_1 _1850_ (.A1(_0796_),
    .A2(_0801_),
    .B1(_1038_),
    .X(_1039_));
 sky130_fd_sc_hd__nand2_1 _1851_ (.A(net54),
    .B(net65),
    .Y(_1040_));
 sky130_fd_sc_hd__xnor2_2 _1852_ (.A(_1039_),
    .B(_1040_),
    .Y(_1041_));
 sky130_fd_sc_hd__inv_2 _1853_ (.A(_1041_),
    .Y(_1042_));
 sky130_fd_sc_hd__xor2_1 _1854_ (.A(_1032_),
    .B(_1035_),
    .X(_1043_));
 sky130_fd_sc_hd__o21ai_2 _1855_ (.A1(_1042_),
    .A2(_1043_),
    .B1(_1036_),
    .Y(_1044_));
 sky130_fd_sc_hd__nand2b_1 _1856_ (.A_N(_1030_),
    .B(_1044_),
    .Y(_1045_));
 sky130_fd_sc_hd__xor2_1 _1857_ (.A(_1030_),
    .B(_1044_),
    .X(_1046_));
 sky130_fd_sc_hd__and4_1 _1858_ (.A(net51),
    .B(net49),
    .C(net69),
    .D(net67),
    .X(_1047_));
 sky130_fd_sc_hd__inv_2 _1859_ (.A(_1047_),
    .Y(_1048_));
 sky130_fd_sc_hd__a22o_1 _1860_ (.A1(net49),
    .A2(net69),
    .B1(net67),
    .B2(net51),
    .X(_1049_));
 sky130_fd_sc_hd__and4_1 _1861_ (.A(net47),
    .B(net70),
    .C(_1048_),
    .D(_1049_),
    .X(_1050_));
 sky130_fd_sc_hd__or2_1 _1862_ (.A(_1047_),
    .B(_1050_),
    .X(_1051_));
 sky130_fd_sc_hd__a31o_1 _1863_ (.A1(net54),
    .A2(\MAC.b[6] ),
    .A3(_1038_),
    .B1(_1037_),
    .X(_1052_));
 sky130_fd_sc_hd__xnor2_1 _1864_ (.A(_1006_),
    .B(_1007_),
    .Y(_1053_));
 sky130_fd_sc_hd__and2_1 _1865_ (.A(_1052_),
    .B(_1053_),
    .X(_1054_));
 sky130_fd_sc_hd__xor2_1 _1866_ (.A(_1052_),
    .B(_1053_),
    .X(_1055_));
 sky130_fd_sc_hd__nor2_1 _1867_ (.A(_1051_),
    .B(_1055_),
    .Y(_1056_));
 sky130_fd_sc_hd__and2_1 _1868_ (.A(_1051_),
    .B(_1055_),
    .X(_1057_));
 sky130_fd_sc_hd__or2_1 _1869_ (.A(_1056_),
    .B(_1057_),
    .X(_1058_));
 sky130_fd_sc_hd__or2_1 _1870_ (.A(_1046_),
    .B(_1058_),
    .X(_1059_));
 sky130_fd_sc_hd__a21o_1 _1871_ (.A1(_1045_),
    .A2(_1059_),
    .B1(_1028_),
    .X(_1060_));
 sky130_fd_sc_hd__nand3_1 _1872_ (.A(_1028_),
    .B(_1045_),
    .C(_1059_),
    .Y(_1061_));
 sky130_fd_sc_hd__o211ai_2 _1873_ (.A1(_1054_),
    .A2(_1057_),
    .B1(_1060_),
    .C1(_1061_),
    .Y(_1062_));
 sky130_fd_sc_hd__a211oi_1 _1874_ (.A1(_1060_),
    .A2(_1062_),
    .B1(_1020_),
    .C1(_1027_),
    .Y(_1063_));
 sky130_fd_sc_hd__o211a_1 _1875_ (.A1(_1020_),
    .A2(_1027_),
    .B1(_1060_),
    .C1(_1062_),
    .X(_1064_));
 sky130_fd_sc_hd__nor2_1 _1876_ (.A(_1063_),
    .B(_1064_),
    .Y(_1065_));
 sky130_fd_sc_hd__and2_1 _1877_ (.A(net72),
    .B(_1065_),
    .X(_1066_));
 sky130_fd_sc_hd__o21ai_1 _1878_ (.A1(_1063_),
    .A2(_1066_),
    .B1(_1026_),
    .Y(_1067_));
 sky130_fd_sc_hd__or3_1 _1879_ (.A(_1026_),
    .B(_1063_),
    .C(_1066_),
    .X(_1068_));
 sky130_fd_sc_hd__nand2_1 _1880_ (.A(_1067_),
    .B(_1068_),
    .Y(_1069_));
 sky130_fd_sc_hd__nor2_1 _1881_ (.A(net72),
    .B(_1065_),
    .Y(_1070_));
 sky130_fd_sc_hd__or2_1 _1882_ (.A(_1066_),
    .B(_1070_),
    .X(_1071_));
 sky130_fd_sc_hd__a211o_1 _1883_ (.A1(_1060_),
    .A2(_1061_),
    .B1(_1054_),
    .C1(_1057_),
    .X(_1072_));
 sky130_fd_sc_hd__nand2_1 _1884_ (.A(_1062_),
    .B(_1072_),
    .Y(_1073_));
 sky130_fd_sc_hd__nand2_1 _1885_ (.A(_1046_),
    .B(_1058_),
    .Y(_1074_));
 sky130_fd_sc_hd__nand2_1 _1886_ (.A(_1059_),
    .B(_1074_),
    .Y(_1075_));
 sky130_fd_sc_hd__xnor2_1 _1887_ (.A(_1041_),
    .B(_1043_),
    .Y(_1076_));
 sky130_fd_sc_hd__a22oi_1 _1888_ (.A1(net56),
    .A2(net64),
    .B1(net62),
    .B2(net58),
    .Y(_1077_));
 sky130_fd_sc_hd__and4_1 _1889_ (.A(net58),
    .B(net56),
    .C(net64),
    .D(net62),
    .X(_0058_));
 sky130_fd_sc_hd__or2_1 _1890_ (.A(_1077_),
    .B(_0058_),
    .X(_0059_));
 sky130_fd_sc_hd__and2_1 _1891_ (.A(net47),
    .B(net76),
    .X(_0060_));
 sky130_fd_sc_hd__nand2_1 _1892_ (.A(net48),
    .B(net76),
    .Y(_0061_));
 sky130_fd_sc_hd__and3_1 _1893_ (.A(net45),
    .B(net73),
    .C(_0061_),
    .X(_0062_));
 sky130_fd_sc_hd__xnor2_1 _1894_ (.A(_1034_),
    .B(_0062_),
    .Y(_0063_));
 sky130_fd_sc_hd__and2b_1 _1895_ (.A_N(_0059_),
    .B(_0063_),
    .X(_0064_));
 sky130_fd_sc_hd__a41o_1 _1896_ (.A1(net46),
    .A2(_0328_),
    .A3(net73),
    .A4(_0060_),
    .B1(_0064_),
    .X(_0065_));
 sky130_fd_sc_hd__a22oi_1 _1897_ (.A1(net47),
    .A2(net70),
    .B1(_1048_),
    .B2(_1049_),
    .Y(_0066_));
 sky130_fd_sc_hd__nor2_1 _1898_ (.A(_1050_),
    .B(_0066_),
    .Y(_0067_));
 sky130_fd_sc_hd__xnor2_1 _1899_ (.A(_0058_),
    .B(_0067_),
    .Y(_0068_));
 sky130_fd_sc_hd__nand3_1 _1900_ (.A(net54),
    .B(net52),
    .C(_0798_),
    .Y(_0069_));
 sky130_fd_sc_hd__a22o_1 _1901_ (.A1(net51),
    .A2(net68),
    .B1(net66),
    .B2(net55),
    .X(_0070_));
 sky130_fd_sc_hd__nand4_1 _1902_ (.A(net49),
    .B(net71),
    .C(_0069_),
    .D(_0070_),
    .Y(_0071_));
 sky130_fd_sc_hd__nand2_1 _1903_ (.A(_0069_),
    .B(_0071_),
    .Y(_0072_));
 sky130_fd_sc_hd__and2b_1 _1904_ (.A_N(_0068_),
    .B(_0072_),
    .X(_0073_));
 sky130_fd_sc_hd__xor2_1 _1905_ (.A(_0068_),
    .B(_0072_),
    .X(_0074_));
 sky130_fd_sc_hd__xnor2_1 _1906_ (.A(_1076_),
    .B(_0065_),
    .Y(_0075_));
 sky130_fd_sc_hd__or2_1 _1907_ (.A(_0074_),
    .B(_0075_),
    .X(_0076_));
 sky130_fd_sc_hd__a21bo_1 _1908_ (.A1(_1076_),
    .A2(_0065_),
    .B1_N(_0076_),
    .X(_0077_));
 sky130_fd_sc_hd__and3_1 _1909_ (.A(_1059_),
    .B(_1074_),
    .C(_0077_),
    .X(_0078_));
 sky130_fd_sc_hd__and2b_1 _1910_ (.A_N(_0077_),
    .B(_1075_),
    .X(_0079_));
 sky130_fd_sc_hd__xnor2_1 _1911_ (.A(_1075_),
    .B(_0077_),
    .Y(_0080_));
 sky130_fd_sc_hd__a21oi_1 _1912_ (.A1(_0058_),
    .A2(_0067_),
    .B1(_0073_),
    .Y(_0081_));
 sky130_fd_sc_hd__o21ba_1 _1913_ (.A1(_0079_),
    .A2(_0081_),
    .B1_N(_0078_),
    .X(_0082_));
 sky130_fd_sc_hd__or2_1 _1914_ (.A(_1073_),
    .B(_0082_),
    .X(_0083_));
 sky130_fd_sc_hd__xnor2_1 _1915_ (.A(_1073_),
    .B(_0082_),
    .Y(_0084_));
 sky130_fd_sc_hd__nand2_1 _1916_ (.A(net42),
    .B(net72),
    .Y(_0085_));
 sky130_fd_sc_hd__or2_1 _1917_ (.A(_0084_),
    .B(_0085_),
    .X(_0086_));
 sky130_fd_sc_hd__a21o_1 _1918_ (.A1(_0083_),
    .A2(_0086_),
    .B1(_1071_),
    .X(_0087_));
 sky130_fd_sc_hd__nand3_1 _1919_ (.A(_1071_),
    .B(_0083_),
    .C(_0086_),
    .Y(_0088_));
 sky130_fd_sc_hd__and2_1 _1920_ (.A(_0087_),
    .B(_0088_),
    .X(_0089_));
 sky130_fd_sc_hd__nand2_1 _1921_ (.A(_0084_),
    .B(_0085_),
    .Y(_0090_));
 sky130_fd_sc_hd__and2_1 _1922_ (.A(_0086_),
    .B(_0090_),
    .X(_0091_));
 sky130_fd_sc_hd__xnor2_1 _1923_ (.A(_0080_),
    .B(_0081_),
    .Y(_0092_));
 sky130_fd_sc_hd__nand2_1 _1924_ (.A(_0074_),
    .B(_0075_),
    .Y(_0093_));
 sky130_fd_sc_hd__xnor2_1 _1925_ (.A(_0059_),
    .B(_0063_),
    .Y(_0094_));
 sky130_fd_sc_hd__nand2_1 _1926_ (.A(net50),
    .B(net73),
    .Y(_0095_));
 sky130_fd_sc_hd__nand2_1 _1927_ (.A(net50),
    .B(net76),
    .Y(_0096_));
 sky130_fd_sc_hd__nor3_1 _1928_ (.A(net46),
    .B(_0061_),
    .C(_0095_),
    .Y(_0097_));
 sky130_fd_sc_hd__nand2_1 _1929_ (.A(net58),
    .B(net64),
    .Y(_0098_));
 sky130_fd_sc_hd__and3_1 _1930_ (.A(net48),
    .B(net74),
    .C(_0096_),
    .X(_0099_));
 sky130_fd_sc_hd__xnor2_1 _1931_ (.A(_1033_),
    .B(_0099_),
    .Y(_0100_));
 sky130_fd_sc_hd__and3_1 _1932_ (.A(net58),
    .B(net64),
    .C(_0100_),
    .X(_0101_));
 sky130_fd_sc_hd__o21a_1 _1933_ (.A1(_0097_),
    .A2(_0101_),
    .B1(_0094_),
    .X(_0102_));
 sky130_fd_sc_hd__a22o_1 _1934_ (.A1(net50),
    .A2(net71),
    .B1(_0069_),
    .B2(_0070_),
    .X(_0103_));
 sky130_fd_sc_hd__and2_1 _1935_ (.A(_0071_),
    .B(_0103_),
    .X(_0104_));
 sky130_fd_sc_hd__and4_1 _1936_ (.A(net56),
    .B(net55),
    .C(net69),
    .D(net67),
    .X(_0105_));
 sky130_fd_sc_hd__inv_2 _1937_ (.A(_0105_),
    .Y(_0106_));
 sky130_fd_sc_hd__a22o_1 _1938_ (.A1(net55),
    .A2(net68),
    .B1(net66),
    .B2(net56),
    .X(_0107_));
 sky130_fd_sc_hd__and4_1 _1939_ (.A(net51),
    .B(net70),
    .C(_0106_),
    .D(_0107_),
    .X(_0108_));
 sky130_fd_sc_hd__o21ai_1 _1940_ (.A1(_0105_),
    .A2(_0108_),
    .B1(_0104_),
    .Y(_0109_));
 sky130_fd_sc_hd__or3_1 _1941_ (.A(_0104_),
    .B(_0105_),
    .C(_0108_),
    .X(_0110_));
 sky130_fd_sc_hd__and2_1 _1942_ (.A(_0109_),
    .B(_0110_),
    .X(_0111_));
 sky130_fd_sc_hd__or3_1 _1943_ (.A(_0094_),
    .B(_0097_),
    .C(_0101_),
    .X(_0112_));
 sky130_fd_sc_hd__and2b_1 _1944_ (.A_N(_0102_),
    .B(_0112_),
    .X(_0113_));
 sky130_fd_sc_hd__and2_1 _1945_ (.A(_0111_),
    .B(_0113_),
    .X(_0114_));
 sky130_fd_sc_hd__o211a_1 _1946_ (.A1(_0102_),
    .A2(_0114_),
    .B1(_0076_),
    .C1(_0093_),
    .X(_0115_));
 sky130_fd_sc_hd__a211oi_1 _1947_ (.A1(_0076_),
    .A2(_0093_),
    .B1(_0102_),
    .C1(_0114_),
    .Y(_0116_));
 sky130_fd_sc_hd__nor3_1 _1948_ (.A(_0109_),
    .B(_0115_),
    .C(_0116_),
    .Y(_0117_));
 sky130_fd_sc_hd__nor2_1 _1949_ (.A(_0115_),
    .B(_0117_),
    .Y(_0118_));
 sky130_fd_sc_hd__and2b_1 _1950_ (.A_N(_0118_),
    .B(_0092_),
    .X(_0119_));
 sky130_fd_sc_hd__xnor2_1 _1951_ (.A(_0092_),
    .B(_0118_),
    .Y(_0120_));
 sky130_fd_sc_hd__nand2_1 _1952_ (.A(net43),
    .B(net72),
    .Y(_0121_));
 sky130_fd_sc_hd__a31o_1 _1953_ (.A1(net43),
    .A2(net72),
    .A3(_0120_),
    .B1(_0119_),
    .X(_0122_));
 sky130_fd_sc_hd__and2_1 _1954_ (.A(_0091_),
    .B(_0122_),
    .X(_0123_));
 sky130_fd_sc_hd__xnor2_1 _1955_ (.A(_0091_),
    .B(_0122_),
    .Y(_0124_));
 sky130_fd_sc_hd__xor2_1 _1956_ (.A(_0120_),
    .B(_0121_),
    .X(_0125_));
 sky130_fd_sc_hd__o21a_1 _1957_ (.A1(_0115_),
    .A2(_0116_),
    .B1(_0109_),
    .X(_0126_));
 sky130_fd_sc_hd__nor2_1 _1958_ (.A(_0117_),
    .B(_0126_),
    .Y(_0127_));
 sky130_fd_sc_hd__xnor2_1 _1959_ (.A(_0111_),
    .B(_0113_),
    .Y(_0128_));
 sky130_fd_sc_hd__xnor2_1 _1960_ (.A(_0098_),
    .B(_0100_),
    .Y(_0129_));
 sky130_fd_sc_hd__nand2_1 _1961_ (.A(net53),
    .B(net75),
    .Y(_0130_));
 sky130_fd_sc_hd__and4_1 _1962_ (.A(net52),
    .B(net50),
    .C(net75),
    .D(net74),
    .X(_0131_));
 sky130_fd_sc_hd__xnor2_1 _1963_ (.A(_0060_),
    .B(_0095_),
    .Y(_0132_));
 sky130_fd_sc_hd__nand2_1 _1964_ (.A(_0061_),
    .B(_0131_),
    .Y(_0133_));
 sky130_fd_sc_hd__and3_1 _1965_ (.A(_0061_),
    .B(_0129_),
    .C(_0131_),
    .X(_0134_));
 sky130_fd_sc_hd__a22oi_1 _1966_ (.A1(net51),
    .A2(net71),
    .B1(_0106_),
    .B2(_0107_),
    .Y(_0135_));
 sky130_fd_sc_hd__nor2_1 _1967_ (.A(_0108_),
    .B(_0135_),
    .Y(_0136_));
 sky130_fd_sc_hd__nor2_1 _1968_ (.A(_0796_),
    .B(_0799_),
    .Y(_0137_));
 sky130_fd_sc_hd__nand2_1 _1969_ (.A(net54),
    .B(net71),
    .Y(_0138_));
 sky130_fd_sc_hd__a22o_1 _1970_ (.A1(net56),
    .A2(net68),
    .B1(net66),
    .B2(net58),
    .X(_0139_));
 sky130_fd_sc_hd__o21a_1 _1971_ (.A1(_0796_),
    .A2(_0799_),
    .B1(_0139_),
    .X(_0140_));
 sky130_fd_sc_hd__a31o_1 _1972_ (.A1(net55),
    .A2(net71),
    .A3(_0139_),
    .B1(_0137_),
    .X(_0141_));
 sky130_fd_sc_hd__nand2_1 _1973_ (.A(_0136_),
    .B(_0141_),
    .Y(_0142_));
 sky130_fd_sc_hd__xor2_1 _1974_ (.A(_0136_),
    .B(_0141_),
    .X(_0143_));
 sky130_fd_sc_hd__xnor2_1 _1975_ (.A(_0129_),
    .B(_0133_),
    .Y(_0144_));
 sky130_fd_sc_hd__a21oi_1 _1976_ (.A1(_0143_),
    .A2(_0144_),
    .B1(_0134_),
    .Y(_0145_));
 sky130_fd_sc_hd__xor2_1 _1977_ (.A(_0128_),
    .B(_0145_),
    .X(_0146_));
 sky130_fd_sc_hd__and3_1 _1978_ (.A(_0136_),
    .B(_0141_),
    .C(_0146_),
    .X(_0147_));
 sky130_fd_sc_hd__o21ba_1 _1979_ (.A1(_0128_),
    .A2(_0145_),
    .B1_N(_0147_),
    .X(_0148_));
 sky130_fd_sc_hd__or3_1 _1980_ (.A(_0117_),
    .B(_0126_),
    .C(_0148_),
    .X(_0149_));
 sky130_fd_sc_hd__nand2_1 _1981_ (.A(net45),
    .B(net72),
    .Y(_0150_));
 sky130_fd_sc_hd__xnor2_1 _1982_ (.A(_0127_),
    .B(_0148_),
    .Y(_0151_));
 sky130_fd_sc_hd__nand2b_1 _1983_ (.A_N(_0150_),
    .B(_0151_),
    .Y(_0152_));
 sky130_fd_sc_hd__a21o_1 _1984_ (.A1(_0149_),
    .A2(_0152_),
    .B1(_0125_),
    .X(_0153_));
 sky130_fd_sc_hd__nand3_1 _1985_ (.A(_0125_),
    .B(_0149_),
    .C(_0152_),
    .Y(_0154_));
 sky130_fd_sc_hd__xnor2_1 _1986_ (.A(_0150_),
    .B(_0151_),
    .Y(_0155_));
 sky130_fd_sc_hd__xnor2_1 _1987_ (.A(_0142_),
    .B(_0146_),
    .Y(_0156_));
 sky130_fd_sc_hd__xnor2_1 _1988_ (.A(_0143_),
    .B(_0144_),
    .Y(_0157_));
 sky130_fd_sc_hd__a22o_1 _1989_ (.A1(net50),
    .A2(net75),
    .B1(net74),
    .B2(net52),
    .X(_0158_));
 sky130_fd_sc_hd__and2b_1 _1990_ (.A_N(_0131_),
    .B(_0158_),
    .X(_0159_));
 sky130_fd_sc_hd__and4_1 _1991_ (.A(net54),
    .B(net52),
    .C(net75),
    .D(net74),
    .X(_0160_));
 sky130_fd_sc_hd__and3b_1 _1992_ (.A_N(_0131_),
    .B(_0158_),
    .C(_0160_),
    .X(_0161_));
 sky130_fd_sc_hd__nand2_1 _1993_ (.A(_0132_),
    .B(_0161_),
    .Y(_0162_));
 sky130_fd_sc_hd__xnor2_1 _1994_ (.A(_0138_),
    .B(_0140_),
    .Y(_0163_));
 sky130_fd_sc_hd__and4_1 _1995_ (.A(net59),
    .B(net57),
    .C(net71),
    .D(net68),
    .X(_0164_));
 sky130_fd_sc_hd__nand2_1 _1996_ (.A(_0163_),
    .B(_0164_),
    .Y(_0165_));
 sky130_fd_sc_hd__xnor2_1 _1997_ (.A(_0163_),
    .B(_0164_),
    .Y(_0166_));
 sky130_fd_sc_hd__or3_1 _1998_ (.A(_0131_),
    .B(_0132_),
    .C(_0161_),
    .X(_0167_));
 sky130_fd_sc_hd__and3_1 _1999_ (.A(_0133_),
    .B(_0162_),
    .C(_0167_),
    .X(_0168_));
 sky130_fd_sc_hd__and2b_1 _2000_ (.A_N(_0166_),
    .B(_0168_),
    .X(_0169_));
 sky130_fd_sc_hd__a21o_1 _2001_ (.A1(_0132_),
    .A2(_0161_),
    .B1(_0169_),
    .X(_0170_));
 sky130_fd_sc_hd__nand2b_1 _2002_ (.A_N(_0157_),
    .B(_0170_),
    .Y(_0171_));
 sky130_fd_sc_hd__xor2_1 _2003_ (.A(_0157_),
    .B(_0170_),
    .X(_0172_));
 sky130_fd_sc_hd__o21a_1 _2004_ (.A1(_0165_),
    .A2(_0172_),
    .B1(_0171_),
    .X(_0173_));
 sky130_fd_sc_hd__and2b_1 _2005_ (.A_N(_0173_),
    .B(_0156_),
    .X(_0174_));
 sky130_fd_sc_hd__nand2_1 _2006_ (.A(net47),
    .B(net72),
    .Y(_0175_));
 sky130_fd_sc_hd__xnor2_1 _2007_ (.A(_0156_),
    .B(_0173_),
    .Y(_0176_));
 sky130_fd_sc_hd__a31o_1 _2008_ (.A1(net47),
    .A2(net72),
    .A3(_0176_),
    .B1(_0174_),
    .X(_0177_));
 sky130_fd_sc_hd__and2_1 _2009_ (.A(_0155_),
    .B(_0177_),
    .X(_0178_));
 sky130_fd_sc_hd__xnor2_1 _2010_ (.A(_0175_),
    .B(_0176_),
    .Y(_0179_));
 sky130_fd_sc_hd__xnor2_1 _2011_ (.A(_0166_),
    .B(_0168_),
    .Y(_0180_));
 sky130_fd_sc_hd__nand2_1 _2012_ (.A(net75),
    .B(_0916_),
    .Y(_0181_));
 sky130_fd_sc_hd__a22o_1 _2013_ (.A1(net57),
    .A2(\MAC.b[3] ),
    .B1(net68),
    .B2(net58),
    .X(_0182_));
 sky130_fd_sc_hd__and2b_1 _2014_ (.A_N(_0164_),
    .B(_0182_),
    .X(_0183_));
 sky130_fd_sc_hd__o21bai_1 _2015_ (.A1(net52),
    .A2(_0181_),
    .B1_N(_0160_),
    .Y(_0184_));
 sky130_fd_sc_hd__xnor2_1 _2016_ (.A(_0159_),
    .B(_0184_),
    .Y(_0185_));
 sky130_fd_sc_hd__or3b_1 _2017_ (.A(_0164_),
    .B(_0185_),
    .C_N(_0182_),
    .X(_0186_));
 sky130_fd_sc_hd__o31ai_2 _2018_ (.A1(net52),
    .A2(_0096_),
    .A3(_0181_),
    .B1(_0186_),
    .Y(_0187_));
 sky130_fd_sc_hd__nand2_1 _2019_ (.A(_0180_),
    .B(_0187_),
    .Y(_0188_));
 sky130_fd_sc_hd__xnor2_1 _2020_ (.A(_0165_),
    .B(_0172_),
    .Y(_0189_));
 sky130_fd_sc_hd__nor2_1 _2021_ (.A(_0188_),
    .B(_0189_),
    .Y(_0190_));
 sky130_fd_sc_hd__nand2_1 _2022_ (.A(net50),
    .B(\MAC.b[2] ),
    .Y(_0191_));
 sky130_fd_sc_hd__nand2_1 _2023_ (.A(_0188_),
    .B(_0189_),
    .Y(_0192_));
 sky130_fd_sc_hd__and2b_1 _2024_ (.A_N(_0190_),
    .B(_0192_),
    .X(_0193_));
 sky130_fd_sc_hd__a31o_1 _2025_ (.A1(net50),
    .A2(net72),
    .A3(_0192_),
    .B1(_0190_),
    .X(_0194_));
 sky130_fd_sc_hd__and2_1 _2026_ (.A(_0179_),
    .B(_0194_),
    .X(_0195_));
 sky130_fd_sc_hd__xnor2_1 _2027_ (.A(_0183_),
    .B(_0185_),
    .Y(_0196_));
 sky130_fd_sc_hd__a22o_1 _2028_ (.A1(net54),
    .A2(net75),
    .B1(net74),
    .B2(net57),
    .X(_0197_));
 sky130_fd_sc_hd__and4b_1 _2029_ (.A_N(_0796_),
    .B(_0800_),
    .C(_0181_),
    .D(_0197_),
    .X(_0198_));
 sky130_fd_sc_hd__and3_1 _2030_ (.A(net54),
    .B(net74),
    .C(_0181_),
    .X(_0199_));
 sky130_fd_sc_hd__xnor2_1 _2031_ (.A(_0130_),
    .B(_0199_),
    .Y(_0200_));
 sky130_fd_sc_hd__and2_1 _2032_ (.A(_0198_),
    .B(_0200_),
    .X(_0201_));
 sky130_fd_sc_hd__xor2_1 _2033_ (.A(_0198_),
    .B(_0200_),
    .X(_0202_));
 sky130_fd_sc_hd__and3_1 _2034_ (.A(net59),
    .B(\MAC.b[3] ),
    .C(_0202_),
    .X(_0203_));
 sky130_fd_sc_hd__a31o_1 _2035_ (.A1(net59),
    .A2(net71),
    .A3(_0202_),
    .B1(_0201_),
    .X(_0204_));
 sky130_fd_sc_hd__nand2_1 _2036_ (.A(_0196_),
    .B(_0204_),
    .Y(_0205_));
 sky130_fd_sc_hd__xor2_1 _2037_ (.A(_0180_),
    .B(_0187_),
    .X(_0206_));
 sky130_fd_sc_hd__xnor2_1 _2038_ (.A(_0205_),
    .B(_0206_),
    .Y(_0207_));
 sky130_fd_sc_hd__and2_1 _2039_ (.A(net52),
    .B(_0207_),
    .X(_0208_));
 sky130_fd_sc_hd__a32oi_1 _2040_ (.A1(_0196_),
    .A2(_0204_),
    .A3(_0206_),
    .B1(_0208_),
    .B2(\MAC.b[2] ),
    .Y(_0209_));
 sky130_fd_sc_hd__xor2_1 _2041_ (.A(_0196_),
    .B(_0204_),
    .X(_0210_));
 sky130_fd_sc_hd__o21ai_1 _2042_ (.A1(net54),
    .A2(_0210_),
    .B1(\MAC.b[2] ),
    .Y(_0211_));
 sky130_fd_sc_hd__nand2_1 _2043_ (.A(\MAC.a[2] ),
    .B(_0210_),
    .Y(_0212_));
 sky130_fd_sc_hd__a21oi_1 _2044_ (.A1(_0181_),
    .A2(_0197_),
    .B1(_0800_),
    .Y(_0213_));
 sky130_fd_sc_hd__a21oi_1 _2045_ (.A1(net59),
    .A2(net71),
    .B1(_0202_),
    .Y(_0214_));
 sky130_fd_sc_hd__a31o_1 _2046_ (.A1(net59),
    .A2(\MAC.a[2] ),
    .A3(net75),
    .B1(net57),
    .X(_0215_));
 sky130_fd_sc_hd__or3b_1 _2047_ (.A(_0203_),
    .B(_0214_),
    .C_N(_0215_),
    .X(_0216_));
 sky130_fd_sc_hd__o31a_1 _2048_ (.A1(_0796_),
    .A2(_0198_),
    .A3(_0213_),
    .B1(_0216_),
    .X(_0217_));
 sky130_fd_sc_hd__a2bb2o_1 _2049_ (.A1_N(net52),
    .A2_N(_0207_),
    .B1(_0212_),
    .B2(_0217_),
    .X(_0218_));
 sky130_fd_sc_hd__o31a_1 _2050_ (.A1(_0208_),
    .A2(_0211_),
    .A3(_0218_),
    .B1(_0209_),
    .X(_0219_));
 sky130_fd_sc_hd__or4_1 _2051_ (.A(_0208_),
    .B(_0209_),
    .C(_0211_),
    .D(_0218_),
    .X(_0220_));
 sky130_fd_sc_hd__xor2_1 _2052_ (.A(_0191_),
    .B(_0193_),
    .X(_0221_));
 sky130_fd_sc_hd__a21oi_1 _2053_ (.A1(_0220_),
    .A2(_0221_),
    .B1(_0219_),
    .Y(_0222_));
 sky130_fd_sc_hd__or2_1 _2054_ (.A(_0179_),
    .B(_0194_),
    .X(_0223_));
 sky130_fd_sc_hd__o221a_1 _2055_ (.A1(_0155_),
    .A2(_0177_),
    .B1(_0195_),
    .B2(_0222_),
    .C1(_0223_),
    .X(_0224_));
 sky130_fd_sc_hd__o211ai_1 _2056_ (.A1(_0178_),
    .A2(_0224_),
    .B1(_0153_),
    .C1(_0154_),
    .Y(_0225_));
 sky130_fd_sc_hd__a21oi_1 _2057_ (.A1(_0153_),
    .A2(_0225_),
    .B1(_0124_),
    .Y(_0226_));
 sky130_fd_sc_hd__o21ai_1 _2058_ (.A1(_0123_),
    .A2(_0226_),
    .B1(_0089_),
    .Y(_0227_));
 sky130_fd_sc_hd__a21o_1 _2059_ (.A1(_0087_),
    .A2(_0227_),
    .B1(_1069_),
    .X(_0228_));
 sky130_fd_sc_hd__a21oi_1 _2060_ (.A1(_1067_),
    .A2(_0228_),
    .B1(_1025_),
    .Y(_0229_));
 sky130_fd_sc_hd__o21a_1 _2061_ (.A1(_1023_),
    .A2(_0229_),
    .B1(_0985_),
    .X(_0230_));
 sky130_fd_sc_hd__o21ai_1 _2062_ (.A1(_0984_),
    .A2(_0230_),
    .B1(_0948_),
    .Y(_0231_));
 sky130_fd_sc_hd__or2_1 _2063_ (.A(_0890_),
    .B(_0907_),
    .X(_0232_));
 sky130_fd_sc_hd__nand2_1 _2064_ (.A(_0908_),
    .B(_0232_),
    .Y(_0233_));
 sky130_fd_sc_hd__a21o_1 _2065_ (.A1(_0946_),
    .A2(_0231_),
    .B1(_0233_),
    .X(_0234_));
 sky130_fd_sc_hd__mux2_1 _2066_ (.A0(_0816_),
    .A1(_0894_),
    .S(_0815_),
    .X(_0235_));
 sky130_fd_sc_hd__a21o_1 _2067_ (.A1(net63),
    .A2(_0813_),
    .B1(_0235_),
    .X(_0236_));
 sky130_fd_sc_hd__o21a_1 _2068_ (.A1(_0897_),
    .A2(_0900_),
    .B1(_0236_),
    .X(_0237_));
 sky130_fd_sc_hd__or3_1 _2069_ (.A(_0897_),
    .B(_0900_),
    .C(_0236_),
    .X(_0238_));
 sky130_fd_sc_hd__and2b_1 _2070_ (.A_N(_0237_),
    .B(_0238_),
    .X(_0239_));
 sky130_fd_sc_hd__nand2_1 _2071_ (.A(_0902_),
    .B(_0905_),
    .Y(_0240_));
 sky130_fd_sc_hd__xnor2_1 _2072_ (.A(_0239_),
    .B(_0240_),
    .Y(_0241_));
 sky130_fd_sc_hd__a21oi_1 _2073_ (.A1(_0908_),
    .A2(_0234_),
    .B1(_0241_),
    .Y(_0242_));
 sky130_fd_sc_hd__o21a_1 _2074_ (.A1(_0237_),
    .A2(_0240_),
    .B1(_0238_),
    .X(_0243_));
 sky130_fd_sc_hd__or2_1 _2075_ (.A(_0242_),
    .B(_0243_),
    .X(_0244_));
 sky130_fd_sc_hd__nor2_1 _2076_ (.A(_0817_),
    .B(_0244_),
    .Y(_0245_));
 sky130_fd_sc_hd__a211o_1 _2077_ (.A1(_0153_),
    .A2(_0154_),
    .B1(_0178_),
    .C1(_0224_),
    .X(_0246_));
 sky130_fd_sc_hd__and2_1 _2078_ (.A(_0225_),
    .B(_0246_),
    .X(_0247_));
 sky130_fd_sc_hd__or4_1 _2079_ (.A(\MAC.a[14] ),
    .B(\MAC.a[13] ),
    .C(net59),
    .D(net57),
    .X(_0248_));
 sky130_fd_sc_hd__or4_1 _2080_ (.A(\MAC.a[10] ),
    .B(\MAC.a[9] ),
    .C(\MAC.a[12] ),
    .D(\MAC.a[11] ),
    .X(_0249_));
 sky130_fd_sc_hd__or4_1 _2081_ (.A(net46),
    .B(net44),
    .C(\MAC.a[8] ),
    .D(\MAC.a[15] ),
    .X(_0250_));
 sky130_fd_sc_hd__or4_1 _2082_ (.A(net54),
    .B(net52),
    .C(net50),
    .D(net48),
    .X(_0251_));
 sky130_fd_sc_hd__or4_1 _2083_ (.A(_0248_),
    .B(_0249_),
    .C(_0250_),
    .D(_0251_),
    .X(_0252_));
 sky130_fd_sc_hd__or4_1 _2084_ (.A(\MAC.b[12] ),
    .B(\MAC.b[11] ),
    .C(\MAC.b[14] ),
    .D(\MAC.b[13] ),
    .X(_0253_));
 sky130_fd_sc_hd__or2_1 _2085_ (.A(\MAC.b[10] ),
    .B(\MAC.b[9] ),
    .X(_0254_));
 sky130_fd_sc_hd__or4_1 _2086_ (.A(net75),
    .B(net74),
    .C(net72),
    .D(\MAC.b[3] ),
    .X(_0255_));
 sky130_fd_sc_hd__or4_1 _2087_ (.A(net65),
    .B(net63),
    .C(net61),
    .D(\MAC.b[15] ),
    .X(_0256_));
 sky130_fd_sc_hd__or4_1 _2088_ (.A(_0874_),
    .B(_0253_),
    .C(_0254_),
    .D(_0256_),
    .X(_0257_));
 sky130_fd_sc_hd__o21a_1 _2089_ (.A1(_0255_),
    .A2(_0257_),
    .B1(_0252_),
    .X(_0258_));
 sky130_fd_sc_hd__inv_2 _2090_ (.A(net30),
    .Y(_0259_));
 sky130_fd_sc_hd__and3_1 _2091_ (.A(_0124_),
    .B(_0153_),
    .C(_0225_),
    .X(_0260_));
 sky130_fd_sc_hd__nor2_1 _2092_ (.A(_0226_),
    .B(_0260_),
    .Y(_0261_));
 sky130_fd_sc_hd__mux2_1 _2093_ (.A0(_0261_),
    .A1(_0247_),
    .S(net19),
    .X(_0262_));
 sky130_fd_sc_hd__nand2_1 _2094_ (.A(net30),
    .B(_0262_),
    .Y(_0263_));
 sky130_fd_sc_hd__a21oi_1 _2095_ (.A1(_0812_),
    .A2(_0263_),
    .B1(_0784_),
    .Y(\MAC.mul.c_mul1[0] ));
 sky130_fd_sc_hd__nand2_1 _2096_ (.A(_0782_),
    .B(_0812_),
    .Y(_0264_));
 sky130_fd_sc_hd__or3_1 _2097_ (.A(_0089_),
    .B(_0123_),
    .C(_0226_),
    .X(_0265_));
 sky130_fd_sc_hd__and2_1 _2098_ (.A(_0227_),
    .B(_0265_),
    .X(_0266_));
 sky130_fd_sc_hd__mux2_1 _2099_ (.A0(_0266_),
    .A1(_0261_),
    .S(net19),
    .X(_0267_));
 sky130_fd_sc_hd__a21o_1 _2100_ (.A1(net30),
    .A2(_0267_),
    .B1(net23),
    .X(_0268_));
 sky130_fd_sc_hd__and2_1 _2101_ (.A(net24),
    .B(_0268_),
    .X(\MAC.mul.c_mul1[1] ));
 sky130_fd_sc_hd__nand3_1 _2102_ (.A(_1069_),
    .B(_0087_),
    .C(_0227_),
    .Y(_0269_));
 sky130_fd_sc_hd__and2_1 _2103_ (.A(_0228_),
    .B(_0269_),
    .X(_0270_));
 sky130_fd_sc_hd__mux2_1 _2104_ (.A0(_0270_),
    .A1(_0266_),
    .S(net19),
    .X(_0271_));
 sky130_fd_sc_hd__a21o_1 _2105_ (.A1(net30),
    .A2(_0271_),
    .B1(net23),
    .X(_0272_));
 sky130_fd_sc_hd__and2_1 _2106_ (.A(net24),
    .B(_0272_),
    .X(\MAC.mul.c_mul1[2] ));
 sky130_fd_sc_hd__and3_1 _2107_ (.A(_1025_),
    .B(_1067_),
    .C(_0228_),
    .X(_0273_));
 sky130_fd_sc_hd__nor2_1 _2108_ (.A(_0229_),
    .B(_0273_),
    .Y(_0274_));
 sky130_fd_sc_hd__mux2_1 _2109_ (.A0(_0274_),
    .A1(_0270_),
    .S(net19),
    .X(_0275_));
 sky130_fd_sc_hd__a21o_1 _2110_ (.A1(net30),
    .A2(_0275_),
    .B1(net23),
    .X(_0276_));
 sky130_fd_sc_hd__and2_1 _2111_ (.A(net24),
    .B(_0276_),
    .X(\MAC.mul.c_mul1[3] ));
 sky130_fd_sc_hd__nor3_1 _2112_ (.A(_0985_),
    .B(_1023_),
    .C(_0229_),
    .Y(_0277_));
 sky130_fd_sc_hd__or2_1 _2113_ (.A(_0230_),
    .B(_0277_),
    .X(_0278_));
 sky130_fd_sc_hd__inv_2 _2114_ (.A(_0278_),
    .Y(_0279_));
 sky130_fd_sc_hd__mux2_1 _2115_ (.A0(_0279_),
    .A1(_0274_),
    .S(net19),
    .X(_0280_));
 sky130_fd_sc_hd__a21o_1 _2116_ (.A1(net30),
    .A2(_0280_),
    .B1(net23),
    .X(_0281_));
 sky130_fd_sc_hd__and2_1 _2117_ (.A(net24),
    .B(_0281_),
    .X(\MAC.mul.c_mul1[4] ));
 sky130_fd_sc_hd__or3_1 _2118_ (.A(_0948_),
    .B(_0984_),
    .C(_0230_),
    .X(_0282_));
 sky130_fd_sc_hd__nand2_1 _2119_ (.A(_0231_),
    .B(_0282_),
    .Y(_0283_));
 sky130_fd_sc_hd__mux2_1 _2120_ (.A0(_0283_),
    .A1(_0278_),
    .S(net19),
    .X(_0284_));
 sky130_fd_sc_hd__nor2_1 _2121_ (.A(_0259_),
    .B(_0284_),
    .Y(_0285_));
 sky130_fd_sc_hd__o21a_1 _2122_ (.A1(net23),
    .A2(_0285_),
    .B1(net24),
    .X(\MAC.mul.c_mul1[5] ));
 sky130_fd_sc_hd__nand2_1 _2123_ (.A(net19),
    .B(_0283_),
    .Y(_0286_));
 sky130_fd_sc_hd__nand3_1 _2124_ (.A(_0946_),
    .B(_0231_),
    .C(_0233_),
    .Y(_0287_));
 sky130_fd_sc_hd__and2_1 _2125_ (.A(_0234_),
    .B(_0287_),
    .X(_0288_));
 sky130_fd_sc_hd__o211a_1 _2126_ (.A1(_0245_),
    .A2(_0288_),
    .B1(_0286_),
    .C1(net30),
    .X(_0289_));
 sky130_fd_sc_hd__o21a_1 _2127_ (.A1(net23),
    .A2(_0289_),
    .B1(net24),
    .X(\MAC.mul.c_mul1[6] ));
 sky130_fd_sc_hd__and3_1 _2128_ (.A(_0908_),
    .B(_0234_),
    .C(_0241_),
    .X(_0290_));
 sky130_fd_sc_hd__nor2_1 _2129_ (.A(_0242_),
    .B(_0290_),
    .Y(_0291_));
 sky130_fd_sc_hd__mux2_1 _2130_ (.A0(_0291_),
    .A1(_0288_),
    .S(net19),
    .X(_0292_));
 sky130_fd_sc_hd__a21o_1 _2131_ (.A1(net30),
    .A2(_0292_),
    .B1(net23),
    .X(_0293_));
 sky130_fd_sc_hd__and2_1 _2132_ (.A(net24),
    .B(_0293_),
    .X(\MAC.mul.c_mul1[7] ));
 sky130_fd_sc_hd__and2_1 _2133_ (.A(_0817_),
    .B(_0244_),
    .X(_0294_));
 sky130_fd_sc_hd__a21o_1 _2134_ (.A1(_0245_),
    .A2(_0291_),
    .B1(_0294_),
    .X(_0295_));
 sky130_fd_sc_hd__a21o_1 _2135_ (.A1(net30),
    .A2(_0295_),
    .B1(net23),
    .X(_0296_));
 sky130_fd_sc_hd__and2_1 _2136_ (.A(net24),
    .B(_0296_),
    .X(\MAC.mul.c_mul1[8] ));
 sky130_fd_sc_hd__nand2_1 _2137_ (.A(_0777_),
    .B(net19),
    .Y(_0297_));
 sky130_fd_sc_hd__or2_1 _2138_ (.A(_0777_),
    .B(net19),
    .X(_0298_));
 sky130_fd_sc_hd__a21o_1 _2139_ (.A1(_0297_),
    .A2(_0298_),
    .B1(_0259_),
    .X(_0299_));
 sky130_fd_sc_hd__a21oi_1 _2140_ (.A1(_0812_),
    .A2(_0299_),
    .B1(_0784_),
    .Y(\MAC.mul.c_mul1[9] ));
 sky130_fd_sc_hd__xor2_1 _2141_ (.A(_0793_),
    .B(_0297_),
    .X(_0300_));
 sky130_fd_sc_hd__a21o_1 _2142_ (.A1(net30),
    .A2(_0300_),
    .B1(net23),
    .X(_0301_));
 sky130_fd_sc_hd__and2_1 _2143_ (.A(net24),
    .B(_0301_),
    .X(\MAC.mul.c_mul1[10] ));
 sky130_fd_sc_hd__o211a_1 _2144_ (.A1(_0817_),
    .A2(_0244_),
    .B1(_0777_),
    .C1(_0793_),
    .X(_0302_));
 sky130_fd_sc_hd__nand2_1 _2145_ (.A(_0792_),
    .B(_0302_),
    .Y(_0303_));
 sky130_fd_sc_hd__o211a_1 _2146_ (.A1(_0792_),
    .A2(_0302_),
    .B1(_0303_),
    .C1(net31),
    .X(_0304_));
 sky130_fd_sc_hd__o21a_1 _2147_ (.A1(net23),
    .A2(_0304_),
    .B1(net24),
    .X(\MAC.mul.c_mul1[11] ));
 sky130_fd_sc_hd__nand3b_1 _2148_ (.A_N(_0788_),
    .B(_0790_),
    .C(_0303_),
    .Y(_0305_));
 sky130_fd_sc_hd__a21bo_1 _2149_ (.A1(_0790_),
    .A2(_0303_),
    .B1_N(_0788_),
    .X(_0306_));
 sky130_fd_sc_hd__a31o_1 _2150_ (.A1(net31),
    .A2(_0305_),
    .A3(_0306_),
    .B1(_0264_),
    .X(_0307_));
 sky130_fd_sc_hd__and2_1 _2151_ (.A(net25),
    .B(_0307_),
    .X(\MAC.mul.c_mul1[12] ));
 sky130_fd_sc_hd__o211a_1 _2152_ (.A1(_0817_),
    .A2(_0244_),
    .B1(_0788_),
    .C1(_0794_),
    .X(_0308_));
 sky130_fd_sc_hd__mux2_1 _2153_ (.A0(_0771_),
    .A1(_0786_),
    .S(_0779_),
    .X(_0309_));
 sky130_fd_sc_hd__and2_1 _2154_ (.A(_0308_),
    .B(_0309_),
    .X(_0310_));
 sky130_fd_sc_hd__o21ai_1 _2155_ (.A1(_0308_),
    .A2(_0309_),
    .B1(net31),
    .Y(_0311_));
 sky130_fd_sc_hd__nor2_1 _2156_ (.A(_0310_),
    .B(_0311_),
    .Y(_0312_));
 sky130_fd_sc_hd__o21a_1 _2157_ (.A1(_0264_),
    .A2(_0312_),
    .B1(net25),
    .X(\MAC.mul.c_mul1[13] ));
 sky130_fd_sc_hd__xor2_1 _2158_ (.A(_0781_),
    .B(_0310_),
    .X(_0313_));
 sky130_fd_sc_hd__a21o_1 _2159_ (.A1(net31),
    .A2(_0313_),
    .B1(_0264_),
    .X(_0314_));
 sky130_fd_sc_hd__and2_1 _2160_ (.A(net25),
    .B(_0314_),
    .X(\MAC.mul.c_mul1[14] ));
 sky130_fd_sc_hd__xor2_1 _2161_ (.A(\MAC.a[15] ),
    .B(\MAC.b[15] ),
    .X(_0315_));
 sky130_fd_sc_hd__a21o_1 _2162_ (.A1(net31),
    .A2(_0315_),
    .B1(_0264_),
    .X(_0316_));
 sky130_fd_sc_hd__o211a_1 _2163_ (.A1(_0782_),
    .A2(_0315_),
    .B1(_0316_),
    .C1(net25),
    .X(\MAC.mul.c_mul1[15] ));
 sky130_fd_sc_hd__mux2_1 _2164_ (.A0(\MAC.add.b1[0] ),
    .A1(\MAC.add.b1[8] ),
    .S(\wrap2.state[0] ),
    .X(_0034_));
 sky130_fd_sc_hd__mux2_1 _2165_ (.A0(\MAC.add.b1[1] ),
    .A1(\MAC.add.b1[9] ),
    .S(\wrap2.state[0] ),
    .X(_0035_));
 sky130_fd_sc_hd__mux2_1 _2166_ (.A0(\MAC.add.b1[2] ),
    .A1(\MAC.add.b1[10] ),
    .S(\wrap2.state[0] ),
    .X(_0036_));
 sky130_fd_sc_hd__mux2_1 _2167_ (.A0(\MAC.add.b1[3] ),
    .A1(\MAC.add.b1[11] ),
    .S(\wrap2.state[0] ),
    .X(_0037_));
 sky130_fd_sc_hd__mux2_1 _2168_ (.A0(\MAC.add.b1[4] ),
    .A1(\MAC.add.b1[12] ),
    .S(\wrap2.state[0] ),
    .X(_0038_));
 sky130_fd_sc_hd__mux2_1 _2169_ (.A0(\MAC.add.b1[5] ),
    .A1(\MAC.add.b1[13] ),
    .S(\wrap2.state[0] ),
    .X(_0039_));
 sky130_fd_sc_hd__mux2_1 _2170_ (.A0(\MAC.add.b1[6] ),
    .A1(\MAC.add.b1[14] ),
    .S(\wrap2.state[0] ),
    .X(_0040_));
 sky130_fd_sc_hd__mux2_1 _2171_ (.A0(\MAC.add.b1[7] ),
    .A1(\MAC.add.b1[15] ),
    .S(\wrap2.state[0] ),
    .X(_0041_));
 sky130_fd_sc_hd__a21o_1 _2172_ (.A1(net35),
    .A2(net2),
    .B1(_0002_),
    .X(_0042_));
 sky130_fd_sc_hd__a21o_1 _2173_ (.A1(net35),
    .A2(net3),
    .B1(_0009_),
    .X(_0043_));
 sky130_fd_sc_hd__a21o_1 _2174_ (.A1(net35),
    .A2(net4),
    .B1(_0010_),
    .X(_0044_));
 sky130_fd_sc_hd__a21o_1 _2175_ (.A1(net36),
    .A2(net5),
    .B1(_0011_),
    .X(_0045_));
 sky130_fd_sc_hd__a21o_1 _2176_ (.A1(net36),
    .A2(net6),
    .B1(_0012_),
    .X(_0046_));
 sky130_fd_sc_hd__a21o_1 _2177_ (.A1(net36),
    .A2(net7),
    .B1(_0013_),
    .X(_0047_));
 sky130_fd_sc_hd__a21o_1 _2178_ (.A1(net36),
    .A2(net8),
    .B1(_0014_),
    .X(_0048_));
 sky130_fd_sc_hd__a21o_1 _2179_ (.A1(net36),
    .A2(net9),
    .B1(_0015_),
    .X(_0049_));
 sky130_fd_sc_hd__a21o_1 _2180_ (.A1(net36),
    .A2(net10),
    .B1(_0016_),
    .X(_0050_));
 sky130_fd_sc_hd__a21o_1 _2181_ (.A1(net35),
    .A2(net11),
    .B1(_0017_),
    .X(_0051_));
 sky130_fd_sc_hd__a21o_1 _2182_ (.A1(net35),
    .A2(net12),
    .B1(_0003_),
    .X(_0052_));
 sky130_fd_sc_hd__a21o_1 _2183_ (.A1(net35),
    .A2(net13),
    .B1(_0004_),
    .X(_0053_));
 sky130_fd_sc_hd__a21o_1 _2184_ (.A1(net35),
    .A2(net14),
    .B1(_0005_),
    .X(_0054_));
 sky130_fd_sc_hd__a21o_1 _2185_ (.A1(net35),
    .A2(net15),
    .B1(_0006_),
    .X(_0055_));
 sky130_fd_sc_hd__a21o_1 _2186_ (.A1(net35),
    .A2(net16),
    .B1(_0007_),
    .X(_0056_));
 sky130_fd_sc_hd__a21o_1 _2187_ (.A1(net35),
    .A2(net17),
    .B1(_0008_),
    .X(_0057_));
 sky130_fd_sc_hd__dfrtp_1 _2188_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0018_),
    .RESET_B(net85),
    .Q(\MAC.b[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2189_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0025_),
    .RESET_B(net85),
    .Q(\MAC.b[1] ));
 sky130_fd_sc_hd__dfrtp_2 _2190_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0026_),
    .RESET_B(net85),
    .Q(\MAC.b[2] ));
 sky130_fd_sc_hd__dfrtp_2 _2191_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0027_),
    .RESET_B(net85),
    .Q(\MAC.b[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2192_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0028_),
    .RESET_B(net85),
    .Q(\MAC.b[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2193_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0029_),
    .RESET_B(net87),
    .Q(\MAC.b[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2194_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0030_),
    .RESET_B(net87),
    .Q(\MAC.b[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2195_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0031_),
    .RESET_B(net87),
    .Q(\MAC.b[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2196_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0032_),
    .RESET_B(net87),
    .Q(\MAC.b[8] ));
 sky130_fd_sc_hd__dfrtp_1 _2197_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0033_),
    .RESET_B(net83),
    .Q(\MAC.b[9] ));
 sky130_fd_sc_hd__dfrtp_1 _2198_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0019_),
    .RESET_B(net83),
    .Q(\MAC.b[10] ));
 sky130_fd_sc_hd__dfrtp_1 _2199_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0020_),
    .RESET_B(net83),
    .Q(\MAC.b[11] ));
 sky130_fd_sc_hd__dfrtp_1 _2200_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0021_),
    .RESET_B(net80),
    .Q(\MAC.b[12] ));
 sky130_fd_sc_hd__dfrtp_2 _2201_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0022_),
    .RESET_B(net80),
    .Q(\MAC.b[13] ));
 sky130_fd_sc_hd__dfrtp_1 _2202_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0023_),
    .RESET_B(net80),
    .Q(\MAC.b[14] ));
 sky130_fd_sc_hd__dfrtp_1 _2203_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0024_),
    .RESET_B(net83),
    .Q(\MAC.b[15] ));
 sky130_fd_sc_hd__dfrtp_4 _2204_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0001_),
    .RESET_B(net78),
    .Q(\wrap2.state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2205_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0002_),
    .RESET_B(net85),
    .Q(\MAC.a[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2206_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0009_),
    .RESET_B(net86),
    .Q(\MAC.a[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2207_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0010_),
    .RESET_B(net85),
    .Q(\MAC.a[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2208_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0011_),
    .RESET_B(net86),
    .Q(\MAC.a[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2209_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0012_),
    .RESET_B(net85),
    .Q(\MAC.a[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2210_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0013_),
    .RESET_B(net86),
    .Q(\MAC.a[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2211_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0014_),
    .RESET_B(net86),
    .Q(\MAC.a[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2212_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0015_),
    .RESET_B(net85),
    .Q(\MAC.a[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2213_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0016_),
    .RESET_B(net83),
    .Q(\MAC.a[8] ));
 sky130_fd_sc_hd__dfrtp_1 _2214_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0017_),
    .RESET_B(net83),
    .Q(\MAC.a[9] ));
 sky130_fd_sc_hd__dfrtp_1 _2215_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0003_),
    .RESET_B(net83),
    .Q(\MAC.a[10] ));
 sky130_fd_sc_hd__dfrtp_1 _2216_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0004_),
    .RESET_B(net84),
    .Q(\MAC.a[11] ));
 sky130_fd_sc_hd__dfrtp_1 _2217_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0005_),
    .RESET_B(net80),
    .Q(\MAC.a[12] ));
 sky130_fd_sc_hd__dfrtp_2 _2218_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0006_),
    .RESET_B(net80),
    .Q(\MAC.a[13] ));
 sky130_fd_sc_hd__dfrtp_1 _2219_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0007_),
    .RESET_B(net80),
    .Q(\MAC.a[14] ));
 sky130_fd_sc_hd__dfrtp_1 _2220_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0008_),
    .RESET_B(net83),
    .Q(\MAC.a[15] ));
 sky130_fd_sc_hd__dfrtp_4 _2221_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0034_),
    .RESET_B(net81),
    .Q(uo_out[0]));
 sky130_fd_sc_hd__dfrtp_4 _2222_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0035_),
    .RESET_B(net81),
    .Q(uo_out[1]));
 sky130_fd_sc_hd__dfrtp_4 _2223_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0036_),
    .RESET_B(net80),
    .Q(uo_out[2]));
 sky130_fd_sc_hd__dfrtp_4 _2224_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0037_),
    .RESET_B(net80),
    .Q(uo_out[3]));
 sky130_fd_sc_hd__dfrtp_4 _2225_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0038_),
    .RESET_B(net81),
    .Q(uo_out[4]));
 sky130_fd_sc_hd__dfrtp_4 _2226_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0039_),
    .RESET_B(net78),
    .Q(uo_out[5]));
 sky130_fd_sc_hd__dfrtp_4 _2227_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0040_),
    .RESET_B(net78),
    .Q(uo_out[6]));
 sky130_fd_sc_hd__dfrtp_4 _2228_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0041_),
    .RESET_B(net79),
    .Q(uo_out[7]));
 sky130_fd_sc_hd__dfrtp_1 _2229_ (.CLK(clknet_3_7__leaf_clk),
    .D(net36),
    .RESET_B(net86),
    .Q(\wrap.state[0] ));
 sky130_fd_sc_hd__dfrtp_2 _2230_ (.CLK(clknet_3_2__leaf_clk),
    .D(\MAC.mul.c_mul1[0] ),
    .RESET_B(net77),
    .Q(\MAC.add.a1[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2231_ (.CLK(clknet_3_2__leaf_clk),
    .D(\MAC.mul.c_mul1[1] ),
    .RESET_B(net77),
    .Q(\MAC.add.a1[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2232_ (.CLK(clknet_3_2__leaf_clk),
    .D(\MAC.mul.c_mul1[2] ),
    .RESET_B(net77),
    .Q(\MAC.add.a1[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2233_ (.CLK(clknet_3_2__leaf_clk),
    .D(\MAC.mul.c_mul1[3] ),
    .RESET_B(net77),
    .Q(\MAC.add.a1[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2234_ (.CLK(clknet_3_2__leaf_clk),
    .D(\MAC.mul.c_mul1[4] ),
    .RESET_B(net77),
    .Q(\MAC.add.a1[4] ));
 sky130_fd_sc_hd__dfrtp_2 _2235_ (.CLK(clknet_3_2__leaf_clk),
    .D(\MAC.mul.c_mul1[5] ),
    .RESET_B(net77),
    .Q(\MAC.add.a1[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2236_ (.CLK(clknet_3_2__leaf_clk),
    .D(\MAC.mul.c_mul1[6] ),
    .RESET_B(net77),
    .Q(\MAC.add.a1[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2237_ (.CLK(clknet_3_2__leaf_clk),
    .D(\MAC.mul.c_mul1[7] ),
    .RESET_B(net77),
    .Q(\MAC.add.a1[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2238_ (.CLK(clknet_3_2__leaf_clk),
    .D(\MAC.mul.c_mul1[8] ),
    .RESET_B(net77),
    .Q(\MAC.add.a1[8] ));
 sky130_fd_sc_hd__dfrtp_4 _2239_ (.CLK(clknet_3_2__leaf_clk),
    .D(\MAC.mul.c_mul1[9] ),
    .RESET_B(net77),
    .Q(\MAC.add.a1[9] ));
 sky130_fd_sc_hd__dfrtp_2 _2240_ (.CLK(clknet_3_3__leaf_clk),
    .D(\MAC.mul.c_mul1[10] ),
    .RESET_B(net82),
    .Q(\MAC.add.a1[10] ));
 sky130_fd_sc_hd__dfrtp_2 _2241_ (.CLK(clknet_3_3__leaf_clk),
    .D(\MAC.mul.c_mul1[11] ),
    .RESET_B(net82),
    .Q(\MAC.add.a1[11] ));
 sky130_fd_sc_hd__dfrtp_4 _2242_ (.CLK(clknet_3_3__leaf_clk),
    .D(\MAC.mul.c_mul1[12] ),
    .RESET_B(net82),
    .Q(\MAC.add.a1[12] ));
 sky130_fd_sc_hd__dfrtp_1 _2243_ (.CLK(clknet_3_3__leaf_clk),
    .D(\MAC.mul.c_mul1[13] ),
    .RESET_B(net82),
    .Q(\MAC.add.a1[13] ));
 sky130_fd_sc_hd__dfrtp_2 _2244_ (.CLK(clknet_3_3__leaf_clk),
    .D(\MAC.mul.c_mul1[14] ),
    .RESET_B(net82),
    .Q(\MAC.add.a1[14] ));
 sky130_fd_sc_hd__dfrtp_1 _2245_ (.CLK(clknet_3_3__leaf_clk),
    .D(\MAC.mul.c_mul1[15] ),
    .RESET_B(net1),
    .Q(\MAC.add.a1[15] ));
 sky130_fd_sc_hd__dfrtp_4 _2246_ (.CLK(clknet_3_0__leaf_clk),
    .D(\MAC.add.c_add[0] ),
    .RESET_B(net78),
    .Q(\MAC.add.b1[0] ));
 sky130_fd_sc_hd__dfrtp_4 _2247_ (.CLK(clknet_3_0__leaf_clk),
    .D(\MAC.add.c_add[1] ),
    .RESET_B(net78),
    .Q(\MAC.add.b1[1] ));
 sky130_fd_sc_hd__dfrtp_4 _2248_ (.CLK(clknet_3_0__leaf_clk),
    .D(\MAC.add.c_add[2] ),
    .RESET_B(net78),
    .Q(\MAC.add.b1[2] ));
 sky130_fd_sc_hd__dfrtp_2 _2249_ (.CLK(clknet_3_0__leaf_clk),
    .D(\MAC.add.c_add[3] ),
    .RESET_B(net82),
    .Q(\MAC.add.b1[3] ));
 sky130_fd_sc_hd__dfrtp_2 _2250_ (.CLK(clknet_3_0__leaf_clk),
    .D(\MAC.add.c_add[4] ),
    .RESET_B(net79),
    .Q(\MAC.add.b1[4] ));
 sky130_fd_sc_hd__dfrtp_4 _2251_ (.CLK(clknet_3_0__leaf_clk),
    .D(\MAC.add.c_add[5] ),
    .RESET_B(net78),
    .Q(\MAC.add.b1[5] ));
 sky130_fd_sc_hd__dfrtp_2 _2252_ (.CLK(clknet_3_0__leaf_clk),
    .D(\MAC.add.c_add[6] ),
    .RESET_B(net78),
    .Q(\MAC.add.b1[6] ));
 sky130_fd_sc_hd__dfrtp_2 _2253_ (.CLK(clknet_3_0__leaf_clk),
    .D(\MAC.add.c_add[7] ),
    .RESET_B(net82),
    .Q(\MAC.add.b1[7] ));
 sky130_fd_sc_hd__dfrtp_4 _2254_ (.CLK(clknet_3_0__leaf_clk),
    .D(\MAC.add.c_add[8] ),
    .RESET_B(net78),
    .Q(\MAC.add.b1[8] ));
 sky130_fd_sc_hd__dfrtp_4 _2255_ (.CLK(clknet_3_3__leaf_clk),
    .D(\MAC.add.c_add[9] ),
    .RESET_B(net82),
    .Q(\MAC.add.b1[9] ));
 sky130_fd_sc_hd__dfrtp_4 _2256_ (.CLK(clknet_3_0__leaf_clk),
    .D(\MAC.add.c_add[10] ),
    .RESET_B(net78),
    .Q(\MAC.add.b1[10] ));
 sky130_fd_sc_hd__dfrtp_4 _2257_ (.CLK(clknet_3_3__leaf_clk),
    .D(\MAC.add.c_add[11] ),
    .RESET_B(net82),
    .Q(\MAC.add.b1[11] ));
 sky130_fd_sc_hd__dfrtp_4 _2258_ (.CLK(clknet_3_0__leaf_clk),
    .D(\MAC.add.c_add[12] ),
    .RESET_B(net79),
    .Q(\MAC.add.b1[12] ));
 sky130_fd_sc_hd__dfrtp_2 _2259_ (.CLK(clknet_3_0__leaf_clk),
    .D(\MAC.add.c_add[13] ),
    .RESET_B(net79),
    .Q(\MAC.add.b1[13] ));
 sky130_fd_sc_hd__dfrtp_2 _2260_ (.CLK(clknet_3_0__leaf_clk),
    .D(\MAC.add.c_add[14] ),
    .RESET_B(net79),
    .Q(\MAC.add.b1[14] ));
 sky130_fd_sc_hd__dfrtp_2 _2261_ (.CLK(clknet_3_3__leaf_clk),
    .D(\MAC.add.c_add[15] ),
    .RESET_B(net1),
    .Q(\MAC.add.b1[15] ));
 sky130_fd_sc_hd__dfrtp_1 _2262_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0042_),
    .RESET_B(net86),
    .Q(\wrap.temp_data[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2263_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0043_),
    .RESET_B(net86),
    .Q(\wrap.temp_data[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2264_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0044_),
    .RESET_B(net86),
    .Q(\wrap.temp_data[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2265_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0045_),
    .RESET_B(net86),
    .Q(\wrap.temp_data[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2266_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0046_),
    .RESET_B(net85),
    .Q(\wrap.temp_data[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2267_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0047_),
    .RESET_B(net84),
    .Q(\wrap.temp_data[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2268_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0048_),
    .RESET_B(net84),
    .Q(\wrap.temp_data[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2269_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0049_),
    .RESET_B(net83),
    .Q(\wrap.temp_data[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2270_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0050_),
    .RESET_B(net83),
    .Q(\wrap.temp_data[8] ));
 sky130_fd_sc_hd__dfrtp_1 _2271_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0051_),
    .RESET_B(net84),
    .Q(\wrap.temp_data[9] ));
 sky130_fd_sc_hd__dfrtp_1 _2272_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0052_),
    .RESET_B(net84),
    .Q(\wrap.temp_data[10] ));
 sky130_fd_sc_hd__dfrtp_1 _2273_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0053_),
    .RESET_B(net84),
    .Q(\wrap.temp_data[11] ));
 sky130_fd_sc_hd__dfrtp_1 _2274_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0054_),
    .RESET_B(net81),
    .Q(\wrap.temp_data[12] ));
 sky130_fd_sc_hd__dfrtp_1 _2275_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0055_),
    .RESET_B(net80),
    .Q(\wrap.temp_data[13] ));
 sky130_fd_sc_hd__dfrtp_1 _2276_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0056_),
    .RESET_B(net81),
    .Q(\wrap.temp_data[14] ));
 sky130_fd_sc_hd__dfrtp_1 _2277_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0057_),
    .RESET_B(net80),
    .Q(\wrap.temp_data[15] ));
 sky130_fd_sc_hd__buf_2 _2278_ (.A(net89),
    .X(uio_oe[0]));
 sky130_fd_sc_hd__buf_2 _2279_ (.A(net90),
    .X(uio_oe[1]));
 sky130_fd_sc_hd__buf_2 _2280_ (.A(net91),
    .X(uio_oe[2]));
 sky130_fd_sc_hd__buf_2 _2281_ (.A(net92),
    .X(uio_oe[3]));
 sky130_fd_sc_hd__buf_2 _2282_ (.A(net93),
    .X(uio_oe[4]));
 sky130_fd_sc_hd__buf_2 _2283_ (.A(net94),
    .X(uio_oe[5]));
 sky130_fd_sc_hd__buf_2 _2284_ (.A(net95),
    .X(uio_oe[6]));
 sky130_fd_sc_hd__buf_2 _2285_ (.A(net96),
    .X(uio_oe[7]));
 sky130_fd_sc_hd__buf_2 _2286_ (.A(net97),
    .X(uio_out[0]));
 sky130_fd_sc_hd__buf_2 _2287_ (.A(net98),
    .X(uio_out[1]));
 sky130_fd_sc_hd__buf_2 _2288_ (.A(net99),
    .X(uio_out[2]));
 sky130_fd_sc_hd__buf_2 _2289_ (.A(net100),
    .X(uio_out[3]));
 sky130_fd_sc_hd__buf_2 _2290_ (.A(net101),
    .X(uio_out[4]));
 sky130_fd_sc_hd__buf_2 _2291_ (.A(net102),
    .X(uio_out[5]));
 sky130_fd_sc_hd__buf_2 _2292_ (.A(net103),
    .X(uio_out[6]));
 sky130_fd_sc_hd__buf_2 _2293_ (.A(net104),
    .X(uio_out[7]));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_617 ();
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(rst_n),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(ui_in[2]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(ui_in[3]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(ui_in[4]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(ui_in[5]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(ui_in[6]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(ui_in[7]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(uio_in[0]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(uio_in[1]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(uio_in[2]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(uio_in[3]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(uio_in[4]),
    .X(net14));
 sky130_fd_sc_hd__buf_1 input15 (.A(uio_in[5]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(uio_in[6]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(uio_in[7]),
    .X(net17));
 sky130_fd_sc_hd__buf_2 fanout18 (.A(_0652_),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_4 fanout19 (.A(_0245_),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 max_cap20 (.A(_0601_),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_4 fanout21 (.A(_0478_),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 fanout22 (.A(_0478_),
    .X(net22));
 sky130_fd_sc_hd__buf_2 fanout23 (.A(_0264_),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 fanout24 (.A(_0783_),
    .X(net24));
 sky130_fd_sc_hd__buf_1 fanout25 (.A(_0783_),
    .X(net25));
 sky130_fd_sc_hd__buf_2 fanout26 (.A(_0391_),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_4 fanout27 (.A(_0351_),
    .X(net27));
 sky130_fd_sc_hd__buf_2 fanout28 (.A(_0351_),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_4 fanout29 (.A(_0350_),
    .X(net29));
 sky130_fd_sc_hd__buf_2 fanout30 (.A(_0258_),
    .X(net30));
 sky130_fd_sc_hd__buf_1 fanout31 (.A(_0258_),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_2 fanout32 (.A(_0365_),
    .X(net32));
 sky130_fd_sc_hd__buf_1 max_cap33 (.A(_0372_),
    .X(net33));
 sky130_fd_sc_hd__buf_2 fanout34 (.A(_0332_),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_4 fanout35 (.A(_0000_),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_2 fanout36 (.A(_0000_),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_2 fanout37 (.A(\wrap.state[0] ),
    .X(net37));
 sky130_fd_sc_hd__buf_1 fanout38 (.A(\wrap.state[0] ),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_2 fanout39 (.A(\wrap.state[0] ),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_2 fanout40 (.A(\wrap.state[0] ),
    .X(net40));
 sky130_fd_sc_hd__buf_2 fanout41 (.A(net42),
    .X(net41));
 sky130_fd_sc_hd__buf_2 fanout42 (.A(\MAC.a[8] ),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_4 fanout43 (.A(net44),
    .X(net43));
 sky130_fd_sc_hd__buf_2 fanout44 (.A(\MAC.a[7] ),
    .X(net44));
 sky130_fd_sc_hd__buf_2 fanout45 (.A(net46),
    .X(net45));
 sky130_fd_sc_hd__buf_2 fanout46 (.A(\MAC.a[6] ),
    .X(net46));
 sky130_fd_sc_hd__buf_2 fanout47 (.A(\MAC.a[5] ),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_2 fanout48 (.A(\MAC.a[5] ),
    .X(net48));
 sky130_fd_sc_hd__buf_2 fanout49 (.A(net50),
    .X(net49));
 sky130_fd_sc_hd__buf_2 fanout50 (.A(\MAC.a[4] ),
    .X(net50));
 sky130_fd_sc_hd__buf_2 fanout51 (.A(net53),
    .X(net51));
 sky130_fd_sc_hd__buf_2 fanout52 (.A(net53),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_2 fanout53 (.A(\MAC.a[3] ),
    .X(net53));
 sky130_fd_sc_hd__buf_2 fanout54 (.A(\MAC.a[2] ),
    .X(net54));
 sky130_fd_sc_hd__buf_2 fanout55 (.A(\MAC.a[2] ),
    .X(net55));
 sky130_fd_sc_hd__buf_2 fanout56 (.A(\MAC.a[1] ),
    .X(net56));
 sky130_fd_sc_hd__buf_2 fanout57 (.A(\MAC.a[1] ),
    .X(net57));
 sky130_fd_sc_hd__buf_2 fanout58 (.A(\MAC.a[0] ),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_2 fanout59 (.A(\MAC.a[0] ),
    .X(net59));
 sky130_fd_sc_hd__buf_2 fanout60 (.A(\MAC.b[8] ),
    .X(net60));
 sky130_fd_sc_hd__buf_1 fanout61 (.A(\MAC.b[8] ),
    .X(net61));
 sky130_fd_sc_hd__buf_2 fanout62 (.A(\MAC.b[7] ),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_2 fanout63 (.A(\MAC.b[7] ),
    .X(net63));
 sky130_fd_sc_hd__buf_2 fanout64 (.A(net65),
    .X(net64));
 sky130_fd_sc_hd__buf_2 fanout65 (.A(\MAC.b[6] ),
    .X(net65));
 sky130_fd_sc_hd__buf_2 fanout66 (.A(net67),
    .X(net66));
 sky130_fd_sc_hd__buf_2 fanout67 (.A(\MAC.b[5] ),
    .X(net67));
 sky130_fd_sc_hd__buf_2 fanout68 (.A(net69),
    .X(net68));
 sky130_fd_sc_hd__buf_2 fanout69 (.A(\MAC.b[4] ),
    .X(net69));
 sky130_fd_sc_hd__buf_2 fanout70 (.A(net71),
    .X(net70));
 sky130_fd_sc_hd__buf_2 fanout71 (.A(\MAC.b[3] ),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_4 fanout72 (.A(\MAC.b[2] ),
    .X(net72));
 sky130_fd_sc_hd__buf_2 fanout73 (.A(\MAC.b[1] ),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_2 fanout74 (.A(\MAC.b[1] ),
    .X(net74));
 sky130_fd_sc_hd__buf_2 fanout75 (.A(net76),
    .X(net75));
 sky130_fd_sc_hd__buf_2 fanout76 (.A(\MAC.b[0] ),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_4 fanout77 (.A(net1),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_4 fanout78 (.A(net88),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_2 fanout79 (.A(net88),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_4 fanout80 (.A(net82),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_2 fanout81 (.A(net88),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_4 fanout82 (.A(net88),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_4 fanout83 (.A(net87),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_2 fanout84 (.A(net87),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_4 fanout85 (.A(net87),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_4 fanout86 (.A(net87),
    .X(net86));
 sky130_fd_sc_hd__buf_2 fanout87 (.A(net88),
    .X(net87));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout88 (.A(net1),
    .X(net88));
 sky130_fd_sc_hd__conb_1 _2278__89 (.LO(net89));
 sky130_fd_sc_hd__conb_1 _2279__90 (.LO(net90));
 sky130_fd_sc_hd__conb_1 _2280__91 (.LO(net91));
 sky130_fd_sc_hd__conb_1 _2281__92 (.LO(net92));
 sky130_fd_sc_hd__conb_1 _2282__93 (.LO(net93));
 sky130_fd_sc_hd__conb_1 _2283__94 (.LO(net94));
 sky130_fd_sc_hd__conb_1 _2284__95 (.LO(net95));
 sky130_fd_sc_hd__conb_1 _2285__96 (.LO(net96));
 sky130_fd_sc_hd__conb_1 _2286__97 (.LO(net97));
 sky130_fd_sc_hd__conb_1 _2287__98 (.LO(net98));
 sky130_fd_sc_hd__conb_1 _2288__99 (.LO(net99));
 sky130_fd_sc_hd__conb_1 _2289__100 (.LO(net100));
 sky130_fd_sc_hd__conb_1 _2290__101 (.LO(net101));
 sky130_fd_sc_hd__conb_1 _2291__102 (.LO(net102));
 sky130_fd_sc_hd__conb_1 _2292__103 (.LO(net103));
 sky130_fd_sc_hd__conb_1 _2293__104 (.LO(net104));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\wrap.temp_data[1] ),
    .X(net105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\wrap.temp_data[6] ),
    .X(net106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\wrap.temp_data[10] ),
    .X(net107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\wrap.temp_data[8] ),
    .X(net108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\wrap.temp_data[12] ),
    .X(net109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\wrap.temp_data[11] ),
    .X(net110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\wrap.temp_data[9] ),
    .X(net111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\wrap.temp_data[0] ),
    .X(net112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\wrap.temp_data[7] ),
    .X(net113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\wrap.temp_data[13] ),
    .X(net114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\wrap.temp_data[14] ),
    .X(net115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\wrap.temp_data[5] ),
    .X(net116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\wrap.temp_data[4] ),
    .X(net117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\wrap.temp_data[3] ),
    .X(net118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\wrap.temp_data[2] ),
    .X(net119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\wrap.temp_data[15] ),
    .X(net120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\wrap2.state[0] ),
    .X(net121));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_87 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_58 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_199 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_334 ();
endmodule
